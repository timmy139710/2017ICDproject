
module imgproc_DW01_dec_0 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15;

  CLKINVX1 U1 ( .A(n15), .Y(n1) );
  OR2X1 U2 ( .A(A[1]), .B(A[0]), .Y(n12) );
  CLKINVX1 U3 ( .A(A[10]), .Y(n2) );
  CLKINVX1 U4 ( .A(A[11]), .Y(n3) );
  AO21X1 U5 ( .A0(n4), .A1(A[9]), .B0(n5), .Y(SUM[9]) );
  OAI2BB1X1 U6 ( .A0N(n6), .A1N(A[8]), .B0(n4), .Y(SUM[8]) );
  OAI2BB1X1 U7 ( .A0N(n7), .A1N(A[7]), .B0(n6), .Y(SUM[7]) );
  OAI2BB1X1 U8 ( .A0N(n8), .A1N(A[6]), .B0(n7), .Y(SUM[6]) );
  OAI2BB1X1 U9 ( .A0N(n9), .A1N(A[5]), .B0(n8), .Y(SUM[5]) );
  OAI2BB1X1 U10 ( .A0N(n10), .A1N(A[4]), .B0(n9), .Y(SUM[4]) );
  OAI2BB1X1 U11 ( .A0N(n11), .A1N(A[3]), .B0(n10), .Y(SUM[3]) );
  OAI2BB1X1 U12 ( .A0N(n12), .A1N(A[2]), .B0(n11), .Y(SUM[2]) );
  OAI2BB1X1 U13 ( .A0N(A[0]), .A1N(A[1]), .B0(n12), .Y(SUM[1]) );
  XOR2X1 U14 ( .A(A[13]), .B(n13), .Y(SUM[13]) );
  NOR2X1 U15 ( .A(A[12]), .B(n14), .Y(n13) );
  XNOR2X1 U16 ( .A(A[12]), .B(n14), .Y(SUM[12]) );
  OAI21XL U17 ( .A0(n1), .A1(n3), .B0(n14), .Y(SUM[11]) );
  NAND2X1 U18 ( .A(n1), .B(n3), .Y(n14) );
  OAI21XL U19 ( .A0(n5), .A1(n2), .B0(n15), .Y(SUM[10]) );
  NAND2X1 U20 ( .A(n5), .B(n2), .Y(n15) );
  NOR2X1 U21 ( .A(n4), .B(A[9]), .Y(n5) );
  OR2X1 U22 ( .A(n6), .B(A[8]), .Y(n4) );
  OR2X1 U23 ( .A(n7), .B(A[7]), .Y(n6) );
  OR2X1 U24 ( .A(n8), .B(A[6]), .Y(n7) );
  OR2X1 U25 ( .A(n9), .B(A[5]), .Y(n8) );
  OR2X1 U26 ( .A(n10), .B(A[4]), .Y(n9) );
  OR2X1 U27 ( .A(n11), .B(A[3]), .Y(n10) );
  OR2X1 U28 ( .A(n12), .B(A[2]), .Y(n11) );
  CLKINVX1 U29 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module imgproc_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module imgproc_DW01_inc_1 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module imgproc_DW01_inc_2 ( A, SUM );
  input [13:0] A;
  output [13:0] SUM;

  wire   [13:2] carry;

  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  XOR2XL U1 ( .A(carry[13]), .B(A[13]), .Y(SUM[13]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module imgproc_DW01_inc_3 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module imgproc_DW01_inc_4 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module imgproc_DW_mult_uns_23 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[3]), .Y(n74) );
  CLKINVX1 U37 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U38 ( .A(a[1]), .Y(n76) );
  CLKINVX1 U39 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U40 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U41 ( .A(a[6]), .Y(n71) );
  CLKINVX1 U42 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U43 ( .A(a[7]), .Y(n70) );
  CLKBUFX3 U44 ( .A(a[0]), .Y(product_3_) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW_mult_uns_22 ( a, product );
  input [7:0] a;
  output [16:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n101, n102, n103, n104, n105, n106, n107, n108;

  ADDFXL U3 ( .A(n19), .B(n102), .CI(n3), .CO(n2), .S(product[15]) );
  ADDFXL U4 ( .A(n21), .B(n20), .CI(n4), .CO(n3), .S(product[14]) );
  ADDFXL U5 ( .A(n23), .B(n22), .CI(n5), .CO(n4), .S(product[13]) );
  ADDFXL U6 ( .A(n25), .B(n24), .CI(n6), .CO(n5), .S(product[12]) );
  ADDFXL U7 ( .A(n26), .B(n29), .CI(n7), .CO(n6), .S(product[11]) );
  ADDFXL U8 ( .A(n30), .B(n34), .CI(n8), .CO(n7), .S(product[10]) );
  ADDFXL U9 ( .A(n36), .B(n35), .CI(n9), .CO(n8), .S(product[9]) );
  ADDFXL U10 ( .A(n37), .B(n41), .CI(n10), .CO(n9), .S(product[8]) );
  ADDFXL U11 ( .A(n43), .B(n42), .CI(n11), .CO(n10), .S(product[7]) );
  ADDFXL U12 ( .A(n44), .B(n47), .CI(n12), .CO(n11), .S(product[6]) );
  ADDFXL U13 ( .A(n48), .B(n49), .CI(n13), .CO(n12), .S(product[5]) );
  ADDFXL U14 ( .A(n50), .B(a[2]), .CI(n14), .CO(n13), .S(product[4]) );
  ADDFXL U15 ( .A(a[3]), .B(a[1]), .CI(n15), .CO(n14), .S(product[3]) );
  ADDHXL U16 ( .A(a[0]), .B(a[2]), .CO(n15), .S(product[2]) );
  ADDHXL U19 ( .A(n101), .B(a[5]), .CO(n19), .S(n20) );
  ADDFXL U20 ( .A(n102), .B(a[7]), .CI(a[4]), .CO(n21), .S(n22) );
  ADDFXL U21 ( .A(a[3]), .B(a[6]), .CI(n27), .CO(n23), .S(n24) );
  ADDFXL U22 ( .A(n31), .B(a[2]), .CI(n28), .CO(n25), .S(n26) );
  ADDHXL U23 ( .A(n101), .B(n103), .CO(n27), .S(n28) );
  ADDFXL U24 ( .A(n33), .B(a[1]), .CI(n32), .CO(n29), .S(n30) );
  ADDHXL U25 ( .A(n102), .B(n104), .CO(n31), .S(n32) );
  CMPR42X1 U26 ( .A(n105), .B(n103), .C(a[0]), .D(a[7]), .ICI(n38), .S(n35), 
        .ICO(n33), .CO(n34) );
  ADDFXL U27 ( .A(n40), .B(a[6]), .CI(n39), .CO(n36), .S(n37) );
  ADDHXL U28 ( .A(n106), .B(n104), .CO(n38), .S(n39) );
  CMPR42X1 U29 ( .A(n107), .B(n105), .C(a[5]), .D(a[7]), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U30 ( .A(a[4]), .B(a[6]), .CI(n46), .CO(n43), .S(n44) );
  ADDFXL U33 ( .A(a[3]), .B(n107), .CI(a[5]), .CO(n47), .S(n48) );
  INVXL U51 ( .A(a[1]), .Y(n107) );
  INVXL U52 ( .A(a[2]), .Y(n106) );
  NAND2XL U53 ( .A(a[0]), .B(a[2]), .Y(n45) );
  CLKINVX1 U54 ( .A(a[4]), .Y(n104) );
  CLKINVX1 U55 ( .A(a[3]), .Y(n105) );
  CLKINVX1 U56 ( .A(a[6]), .Y(n102) );
  CLKINVX1 U57 ( .A(a[5]), .Y(n103) );
  CLKINVX1 U58 ( .A(a[7]), .Y(n101) );
  CLKBUFX3 U59 ( .A(a[1]), .Y(product[1]) );
  CLKBUFX3 U60 ( .A(a[0]), .Y(product[0]) );
  XOR2X1 U61 ( .A(n102), .B(n108), .Y(product[16]) );
  XOR2X1 U62 ( .A(n2), .B(a[7]), .Y(n108) );
  XOR2X1 U63 ( .A(a[4]), .B(a[0]), .Y(n50) );
  NAND2X1 U64 ( .A(a[0]), .B(n104), .Y(n49) );
  XOR2X1 U65 ( .A(n106), .B(a[0]), .Y(n46) );
endmodule


module imgproc_DW_mult_uns_21 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U37 ( .A(a[1]), .Y(n76) );
  CLKINVX1 U38 ( .A(a[3]), .Y(n74) );
  CLKINVX1 U39 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U40 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U41 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U42 ( .A(a[6]), .Y(n71) );
  CLKINVX1 U43 ( .A(a[7]), .Y(n70) );
  CLKBUFX3 U44 ( .A(a[0]), .Y(product_3_) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW_mult_uns_19 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U37 ( .A(a[1]), .Y(n76) );
  CLKINVX1 U38 ( .A(a[3]), .Y(n74) );
  CLKINVX1 U39 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U40 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U41 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U42 ( .A(a[7]), .Y(n70) );
  CLKINVX1 U43 ( .A(a[6]), .Y(n71) );
  CLKBUFX3 U44 ( .A(a[0]), .Y(product_3_) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW_mult_uns_17 ( a, product );
  input [7:0] a;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n89, n90,
         n91, n92, n93, n94, n95, n96, n97;

  ADDFXL U3 ( .A(n90), .B(a[5]), .CI(n3), .CO(n2), .S(product[18]) );
  ADDFXL U4 ( .A(n20), .B(n91), .CI(n4), .CO(n3), .S(product[17]) );
  ADDFXL U5 ( .A(n21), .B(n22), .CI(n5), .CO(n4), .S(product[16]) );
  ADDFXL U6 ( .A(n23), .B(n24), .CI(n6), .CO(n5), .S(product[15]) );
  ADDFXL U7 ( .A(n26), .B(n25), .CI(n7), .CO(n6), .S(product[14]) );
  ADDFXL U8 ( .A(n27), .B(n28), .CI(n8), .CO(n7), .S(product[13]) );
  ADDFXL U9 ( .A(n29), .B(n30), .CI(n9), .CO(n8), .S(product[12]) );
  ADDFXL U10 ( .A(n31), .B(n32), .CI(n10), .CO(n9), .S(product[11]) );
  ADDFXL U11 ( .A(n33), .B(a[4]), .CI(n11), .CO(n10), .S(product[10]) );
  ADDFXL U12 ( .A(a[3]), .B(a[0]), .CI(n12), .CO(n11), .S(product[9]) );
  ADDHXL U13 ( .A(a[2]), .B(n13), .CO(n12), .S(product[8]) );
  ADDFXL U14 ( .A(a[7]), .B(a[1]), .CI(n14), .CO(n13), .S(product[7]) );
  ADDHXL U15 ( .A(a[0]), .B(a[6]), .CO(n14), .S(product[6]) );
  ADDHXL U19 ( .A(n89), .B(a[4]), .CO(n20), .S(n21) );
  ADDHXL U20 ( .A(n90), .B(a[3]), .CO(n22), .S(n23) );
  ADDHXL U21 ( .A(n91), .B(a[2]), .CO(n24), .S(n25) );
  ADDFXL U22 ( .A(a[1]), .B(n92), .CI(a[7]), .CO(n26), .S(n27) );
  ADDFXL U23 ( .A(a[0]), .B(n93), .CI(a[6]), .CO(n28), .S(n29) );
  ADDHXL U24 ( .A(n94), .B(a[5]), .CO(n30), .S(n31) );
  ADDHXL U25 ( .A(n96), .B(n95), .CO(n32), .S(n33) );
  CLKINVX1 U41 ( .A(a[1]), .Y(n95) );
  CLKINVX1 U42 ( .A(a[0]), .Y(n96) );
  CLKINVX1 U43 ( .A(a[2]), .Y(n94) );
  CLKINVX1 U44 ( .A(a[3]), .Y(n93) );
  CLKINVX1 U45 ( .A(a[4]), .Y(n92) );
  CLKINVX1 U46 ( .A(a[6]), .Y(n90) );
  CLKINVX1 U47 ( .A(a[5]), .Y(n91) );
  CLKINVX1 U48 ( .A(a[7]), .Y(n89) );
  CLKBUFX3 U49 ( .A(a[5]), .Y(product[5]) );
  CLKBUFX3 U50 ( .A(a[4]), .Y(product[4]) );
  CLKBUFX3 U51 ( .A(a[3]), .Y(product[3]) );
  CLKBUFX3 U52 ( .A(a[2]), .Y(product[2]) );
  CLKBUFX3 U53 ( .A(a[1]), .Y(product[1]) );
  CLKBUFX3 U54 ( .A(a[0]), .Y(product[0]) );
  XOR2X1 U55 ( .A(n90), .B(n97), .Y(product[19]) );
  XOR2X1 U56 ( .A(n2), .B(a[7]), .Y(n97) );
endmodule


module imgproc_DW_mult_uns_15 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U37 ( .A(a[1]), .Y(n76) );
  CLKINVX1 U38 ( .A(a[3]), .Y(n74) );
  CLKINVX1 U39 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U40 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U41 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U42 ( .A(a[7]), .Y(n70) );
  CLKINVX1 U43 ( .A(a[6]), .Y(n71) );
  CLKBUFX3 U44 ( .A(a[0]), .Y(product_3_) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW_mult_uns_14 ( a, product );
  input [7:0] a;
  output [16:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n101, n102, n103, n104, n105, n106, n107, n108;

  ADDFXL U3 ( .A(n19), .B(n102), .CI(n3), .CO(n2), .S(product[15]) );
  ADDFXL U4 ( .A(n21), .B(n20), .CI(n4), .CO(n3), .S(product[14]) );
  ADDFXL U5 ( .A(n23), .B(n22), .CI(n5), .CO(n4), .S(product[13]) );
  ADDFXL U6 ( .A(n25), .B(n24), .CI(n6), .CO(n5), .S(product[12]) );
  ADDFXL U7 ( .A(n26), .B(n29), .CI(n7), .CO(n6), .S(product[11]) );
  ADDFXL U8 ( .A(n30), .B(n34), .CI(n8), .CO(n7), .S(product[10]) );
  ADDFXL U9 ( .A(n36), .B(n35), .CI(n9), .CO(n8), .S(product[9]) );
  ADDFXL U10 ( .A(n37), .B(n41), .CI(n10), .CO(n9), .S(product[8]) );
  ADDFXL U11 ( .A(n43), .B(n42), .CI(n11), .CO(n10), .S(product[7]) );
  ADDFXL U12 ( .A(n44), .B(n47), .CI(n12), .CO(n11), .S(product[6]) );
  ADDFXL U13 ( .A(n48), .B(n49), .CI(n13), .CO(n12), .S(product[5]) );
  ADDFXL U14 ( .A(n50), .B(a[2]), .CI(n14), .CO(n13), .S(product[4]) );
  ADDFXL U15 ( .A(a[3]), .B(a[1]), .CI(n15), .CO(n14), .S(product[3]) );
  ADDHXL U16 ( .A(a[0]), .B(a[2]), .CO(n15), .S(product[2]) );
  ADDHXL U19 ( .A(n101), .B(a[5]), .CO(n19), .S(n20) );
  ADDFXL U20 ( .A(n102), .B(a[7]), .CI(a[4]), .CO(n21), .S(n22) );
  ADDFXL U21 ( .A(a[3]), .B(a[6]), .CI(n27), .CO(n23), .S(n24) );
  ADDFXL U22 ( .A(n31), .B(a[2]), .CI(n28), .CO(n25), .S(n26) );
  ADDHXL U23 ( .A(n101), .B(n103), .CO(n27), .S(n28) );
  ADDFXL U24 ( .A(n33), .B(a[1]), .CI(n32), .CO(n29), .S(n30) );
  ADDHXL U25 ( .A(n102), .B(n104), .CO(n31), .S(n32) );
  CMPR42X1 U26 ( .A(n105), .B(n103), .C(a[0]), .D(a[7]), .ICI(n38), .S(n35), 
        .ICO(n33), .CO(n34) );
  ADDFXL U27 ( .A(n40), .B(a[6]), .CI(n39), .CO(n36), .S(n37) );
  ADDHXL U28 ( .A(n106), .B(n104), .CO(n38), .S(n39) );
  CMPR42X1 U29 ( .A(n107), .B(n105), .C(a[5]), .D(a[7]), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U30 ( .A(a[4]), .B(a[6]), .CI(n46), .CO(n43), .S(n44) );
  ADDFXL U33 ( .A(a[3]), .B(n107), .CI(a[5]), .CO(n47), .S(n48) );
  INVXL U51 ( .A(a[1]), .Y(n107) );
  INVXL U52 ( .A(a[2]), .Y(n106) );
  NAND2XL U53 ( .A(a[0]), .B(a[2]), .Y(n45) );
  CLKINVX1 U54 ( .A(a[4]), .Y(n104) );
  CLKINVX1 U55 ( .A(a[3]), .Y(n105) );
  CLKINVX1 U56 ( .A(a[6]), .Y(n102) );
  CLKINVX1 U57 ( .A(a[5]), .Y(n103) );
  CLKINVX1 U58 ( .A(a[7]), .Y(n101) );
  CLKBUFX3 U59 ( .A(a[1]), .Y(product[1]) );
  CLKBUFX3 U60 ( .A(a[0]), .Y(product[0]) );
  XOR2X1 U61 ( .A(n102), .B(n108), .Y(product[16]) );
  XOR2X1 U62 ( .A(n2), .B(a[7]), .Y(n108) );
  XOR2X1 U63 ( .A(a[4]), .B(a[0]), .Y(n50) );
  NAND2X1 U64 ( .A(a[0]), .B(n104), .Y(n49) );
  XOR2X1 U65 ( .A(n106), .B(a[0]), .Y(n46) );
endmodule


module imgproc_DW_mult_uns_13 ( a, product );
  input [7:0] a;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n89, n90,
         n91, n92, n93, n94, n95, n96, n97;

  ADDFXL U3 ( .A(n90), .B(a[5]), .CI(n3), .CO(n2), .S(product[18]) );
  ADDFXL U4 ( .A(n20), .B(n91), .CI(n4), .CO(n3), .S(product[17]) );
  ADDFXL U5 ( .A(n21), .B(n22), .CI(n5), .CO(n4), .S(product[16]) );
  ADDFXL U6 ( .A(n23), .B(n24), .CI(n6), .CO(n5), .S(product[15]) );
  ADDFXL U7 ( .A(n26), .B(n25), .CI(n7), .CO(n6), .S(product[14]) );
  ADDFXL U8 ( .A(n27), .B(n28), .CI(n8), .CO(n7), .S(product[13]) );
  ADDFXL U9 ( .A(n29), .B(n30), .CI(n9), .CO(n8), .S(product[12]) );
  ADDFXL U10 ( .A(n31), .B(n32), .CI(n10), .CO(n9), .S(product[11]) );
  ADDFXL U11 ( .A(n33), .B(a[4]), .CI(n11), .CO(n10), .S(product[10]) );
  ADDFXL U12 ( .A(a[3]), .B(a[0]), .CI(n12), .CO(n11), .S(product[9]) );
  ADDHXL U13 ( .A(a[2]), .B(n13), .CO(n12), .S(product[8]) );
  ADDFXL U14 ( .A(a[7]), .B(a[1]), .CI(n14), .CO(n13), .S(product[7]) );
  ADDHXL U15 ( .A(a[0]), .B(a[6]), .CO(n14), .S(product[6]) );
  ADDHXL U19 ( .A(n89), .B(a[4]), .CO(n20), .S(n21) );
  ADDHXL U20 ( .A(n90), .B(a[3]), .CO(n22), .S(n23) );
  ADDHXL U21 ( .A(n91), .B(a[2]), .CO(n24), .S(n25) );
  ADDFXL U22 ( .A(a[1]), .B(n92), .CI(a[7]), .CO(n26), .S(n27) );
  ADDFXL U23 ( .A(a[0]), .B(n93), .CI(a[6]), .CO(n28), .S(n29) );
  ADDHXL U24 ( .A(n94), .B(a[5]), .CO(n30), .S(n31) );
  ADDHXL U25 ( .A(n96), .B(n95), .CO(n32), .S(n33) );
  CLKINVX1 U41 ( .A(a[1]), .Y(n95) );
  CLKINVX1 U42 ( .A(a[0]), .Y(n96) );
  CLKINVX1 U43 ( .A(a[2]), .Y(n94) );
  CLKINVX1 U44 ( .A(a[3]), .Y(n93) );
  CLKINVX1 U45 ( .A(a[4]), .Y(n92) );
  CLKINVX1 U46 ( .A(a[6]), .Y(n90) );
  CLKINVX1 U47 ( .A(a[5]), .Y(n91) );
  CLKINVX1 U48 ( .A(a[7]), .Y(n89) );
  CLKBUFX3 U49 ( .A(a[5]), .Y(product[5]) );
  CLKBUFX3 U50 ( .A(a[4]), .Y(product[4]) );
  CLKBUFX3 U51 ( .A(a[3]), .Y(product[3]) );
  CLKBUFX3 U52 ( .A(a[2]), .Y(product[2]) );
  CLKBUFX3 U53 ( .A(a[1]), .Y(product[1]) );
  CLKBUFX3 U54 ( .A(a[0]), .Y(product[0]) );
  XOR2X1 U55 ( .A(n90), .B(n97), .Y(product[19]) );
  XOR2X1 U56 ( .A(n2), .B(a[7]), .Y(n97) );
endmodule


module imgproc_DW_mult_uns_12 ( a, product_20_, product_19_, product_18_, 
        product_17_, product_16_, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_20_, product_19_, product_18_, product_17_, product_16_,
         product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n111, n112, n113, n114, n115, n116,
         n117, n118;

  ADDFXL U3 ( .A(n20), .B(n112), .CI(n3), .CO(n2), .S(product_19_) );
  ADDFXL U4 ( .A(n22), .B(n21), .CI(n4), .CO(n3), .S(product_18_) );
  ADDFXL U5 ( .A(n24), .B(n23), .CI(n5), .CO(n4), .S(product_17_) );
  ADDFXL U6 ( .A(n26), .B(n25), .CI(n6), .CO(n5), .S(product_16_) );
  ADDFXL U7 ( .A(n27), .B(n30), .CI(n7), .CO(n6), .S(product_15_) );
  ADDFXL U8 ( .A(n31), .B(n34), .CI(n8), .CO(n7), .S(product_14_) );
  ADDFXL U9 ( .A(n35), .B(n38), .CI(n9), .CO(n8), .S(product_13_) );
  ADDFXL U10 ( .A(n39), .B(n42), .CI(n10), .CO(n9), .S(product_12_) );
  ADDFXL U11 ( .A(n43), .B(n46), .CI(n11), .CO(n10), .S(product_11_) );
  ADDFXL U12 ( .A(n47), .B(n50), .CI(n12), .CO(n11), .S(product_10_) );
  ADDFXL U13 ( .A(n51), .B(n52), .CI(n13), .CO(n12), .S(product_9_) );
  ADDFXL U14 ( .A(n53), .B(a[0]), .CI(n14), .CO(n13), .S(product_8_) );
  ADDFXL U15 ( .A(a[4]), .B(n116), .CI(n15), .CO(n14), .S(product_7_) );
  ADDFXL U16 ( .A(a[3]), .B(n117), .CI(n16), .CO(n15), .S(product_6_) );
  ADDHXL U22 ( .A(n111), .B(a[5]), .CO(n20), .S(n21) );
  ADDFXL U23 ( .A(n112), .B(a[7]), .CI(a[4]), .CO(n22), .S(n23) );
  ADDFXL U24 ( .A(a[3]), .B(a[6]), .CI(n28), .CO(n24), .S(n25) );
  ADDFXL U25 ( .A(n32), .B(a[2]), .CI(n29), .CO(n26), .S(n27) );
  ADDFXL U28 ( .A(n36), .B(a[1]), .CI(n33), .CO(n30), .S(n31) );
  ADDFXL U31 ( .A(n40), .B(a[0]), .CI(n37), .CO(n34), .S(n35) );
  ADDFXL U34 ( .A(n44), .B(a[4]), .CI(n41), .CO(n38), .S(n39) );
  ADDHXL U35 ( .A(n111), .B(n116), .CO(n40), .S(n41) );
  ADDFXL U36 ( .A(n48), .B(a[3]), .CI(n45), .CO(n42), .S(n43) );
  ADDHXL U37 ( .A(n112), .B(n117), .CO(n44), .S(n45) );
  ADDFXL U38 ( .A(a[2]), .B(a[7]), .CI(n49), .CO(n46), .S(n47) );
  ADDFXL U41 ( .A(a[1]), .B(n114), .CI(a[6]), .CO(n50), .S(n51) );
  ADDHXL U42 ( .A(n115), .B(a[5]), .CO(n52), .S(n53) );
  CLKBUFX2 U59 ( .A(a[0]), .Y(product_3_) );
  NAND2XL U60 ( .A(a[5]), .B(n111), .Y(n28) );
  XNOR2XL U61 ( .A(n111), .B(a[5]), .Y(n29) );
  INVXL U62 ( .A(a[5]), .Y(n113) );
  NAND2XL U63 ( .A(a[5]), .B(a[0]), .Y(n48) );
  XNOR2XL U64 ( .A(a[0]), .B(a[5]), .Y(n49) );
  CLKINVX1 U65 ( .A(a[2]), .Y(n116) );
  CLKINVX1 U66 ( .A(a[1]), .Y(n117) );
  CLKINVX1 U67 ( .A(a[3]), .Y(n115) );
  CLKINVX1 U68 ( .A(a[4]), .Y(n114) );
  CLKINVX1 U69 ( .A(a[7]), .Y(n111) );
  CLKINVX1 U70 ( .A(a[6]), .Y(n112) );
  CLKBUFX3 U71 ( .A(a[1]), .Y(product_4_) );
  XNOR2X1 U72 ( .A(n116), .B(a[0]), .Y(product_5_) );
  XNOR2X1 U73 ( .A(a[6]), .B(n118), .Y(product_20_) );
  XNOR2X1 U74 ( .A(n2), .B(n111), .Y(n118) );
  XNOR2X1 U75 ( .A(n113), .B(a[3]), .Y(n37) );
  NAND2X1 U76 ( .A(a[3]), .B(n113), .Y(n36) );
  XNOR2X1 U77 ( .A(n112), .B(a[4]), .Y(n33) );
  NAND2X1 U78 ( .A(a[4]), .B(n112), .Y(n32) );
  NAND2X1 U79 ( .A(a[0]), .B(n116), .Y(n16) );
endmodule


module imgproc_DW_mult_uns_11 ( a, product );
  input [7:0] a;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n89, n90,
         n91, n92, n93, n94, n95, n96, n97;

  ADDFXL U3 ( .A(n90), .B(a[5]), .CI(n3), .CO(n2), .S(product[18]) );
  ADDFXL U4 ( .A(n20), .B(n91), .CI(n4), .CO(n3), .S(product[17]) );
  ADDFXL U5 ( .A(n21), .B(n22), .CI(n5), .CO(n4), .S(product[16]) );
  ADDFXL U6 ( .A(n23), .B(n24), .CI(n6), .CO(n5), .S(product[15]) );
  ADDFXL U7 ( .A(n26), .B(n25), .CI(n7), .CO(n6), .S(product[14]) );
  ADDFXL U8 ( .A(n27), .B(n28), .CI(n8), .CO(n7), .S(product[13]) );
  ADDFXL U9 ( .A(n29), .B(n30), .CI(n9), .CO(n8), .S(product[12]) );
  ADDFXL U10 ( .A(n31), .B(n32), .CI(n10), .CO(n9), .S(product[11]) );
  ADDFXL U11 ( .A(n33), .B(a[4]), .CI(n11), .CO(n10), .S(product[10]) );
  ADDFXL U12 ( .A(a[3]), .B(a[0]), .CI(n12), .CO(n11), .S(product[9]) );
  ADDHXL U13 ( .A(a[2]), .B(n13), .CO(n12), .S(product[8]) );
  ADDFXL U14 ( .A(a[7]), .B(a[1]), .CI(n14), .CO(n13), .S(product[7]) );
  ADDHXL U15 ( .A(a[0]), .B(a[6]), .CO(n14), .S(product[6]) );
  ADDHXL U19 ( .A(n89), .B(a[4]), .CO(n20), .S(n21) );
  ADDHXL U20 ( .A(n90), .B(a[3]), .CO(n22), .S(n23) );
  ADDHXL U21 ( .A(n91), .B(a[2]), .CO(n24), .S(n25) );
  ADDFXL U22 ( .A(a[1]), .B(n92), .CI(a[7]), .CO(n26), .S(n27) );
  ADDFXL U23 ( .A(a[0]), .B(n93), .CI(a[6]), .CO(n28), .S(n29) );
  ADDHXL U24 ( .A(n94), .B(a[5]), .CO(n30), .S(n31) );
  ADDHXL U25 ( .A(n96), .B(n95), .CO(n32), .S(n33) );
  CLKBUFX3 U41 ( .A(a[1]), .Y(product[1]) );
  CLKBUFX3 U42 ( .A(a[2]), .Y(product[2]) );
  CLKBUFX3 U43 ( .A(a[3]), .Y(product[3]) );
  CLKBUFX3 U44 ( .A(a[0]), .Y(product[0]) );
  CLKBUFX3 U45 ( .A(a[4]), .Y(product[4]) );
  CLKINVX1 U46 ( .A(a[1]), .Y(n95) );
  CLKINVX1 U47 ( .A(a[0]), .Y(n96) );
  CLKINVX1 U48 ( .A(a[2]), .Y(n94) );
  CLKINVX1 U49 ( .A(a[3]), .Y(n93) );
  CLKINVX1 U50 ( .A(a[4]), .Y(n92) );
  CLKINVX1 U51 ( .A(a[6]), .Y(n90) );
  CLKINVX1 U52 ( .A(a[5]), .Y(n91) );
  CLKINVX1 U53 ( .A(a[7]), .Y(n89) );
  CLKBUFX3 U54 ( .A(a[5]), .Y(product[5]) );
  XOR2X1 U55 ( .A(n90), .B(n97), .Y(product[19]) );
  XOR2X1 U56 ( .A(n2), .B(a[7]), .Y(n97) );
endmodule


module imgproc_DW_mult_uns_10 ( a, product );
  input [7:0] a;
  output [16:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n99, n100, n103, n104, n105, n106, n107, n108, n109,
         n110;

  ADDFXL U3 ( .A(n19), .B(n104), .CI(n3), .CO(n2), .S(product[15]) );
  ADDFXL U4 ( .A(n21), .B(n20), .CI(n4), .CO(n3), .S(product[14]) );
  ADDFXL U5 ( .A(n23), .B(n22), .CI(n5), .CO(n4), .S(product[13]) );
  ADDFXL U6 ( .A(n25), .B(n24), .CI(n6), .CO(n5), .S(product[12]) );
  ADDFXL U7 ( .A(n26), .B(n29), .CI(n7), .CO(n6), .S(product[11]) );
  ADDFXL U8 ( .A(n30), .B(n34), .CI(n8), .CO(n7), .S(product[10]) );
  ADDFXL U9 ( .A(n36), .B(n35), .CI(n9), .CO(n8), .S(product[9]) );
  ADDFXL U10 ( .A(n37), .B(n41), .CI(n10), .CO(n9), .S(product[8]) );
  ADDFXL U11 ( .A(n43), .B(n42), .CI(n11), .CO(n10), .S(product[7]) );
  ADDFXL U12 ( .A(n44), .B(n47), .CI(n12), .CO(n11), .S(product[6]) );
  ADDFXL U13 ( .A(n48), .B(n49), .CI(n13), .CO(n12), .S(product[5]) );
  ADDFXL U14 ( .A(n50), .B(n100), .CI(n14), .CO(n13), .S(product[4]) );
  ADDFXL U15 ( .A(a[3]), .B(n99), .CI(n15), .CO(n14), .S(product[3]) );
  ADDHXL U16 ( .A(a[0]), .B(n100), .CO(n15), .S(product[2]) );
  ADDHXL U19 ( .A(n103), .B(a[5]), .CO(n19), .S(n20) );
  ADDFXL U20 ( .A(n104), .B(a[7]), .CI(a[4]), .CO(n21), .S(n22) );
  ADDFXL U21 ( .A(a[3]), .B(a[6]), .CI(n27), .CO(n23), .S(n24) );
  ADDFXL U22 ( .A(n31), .B(n100), .CI(n28), .CO(n25), .S(n26) );
  ADDHXL U23 ( .A(n103), .B(n105), .CO(n27), .S(n28) );
  ADDFXL U24 ( .A(n33), .B(n99), .CI(n32), .CO(n29), .S(n30) );
  ADDHXL U25 ( .A(n104), .B(n106), .CO(n31), .S(n32) );
  CMPR42X1 U26 ( .A(n107), .B(n105), .C(a[0]), .D(a[7]), .ICI(n38), .S(n35), 
        .ICO(n33), .CO(n34) );
  ADDFXL U27 ( .A(n40), .B(a[6]), .CI(n39), .CO(n36), .S(n37) );
  ADDHXL U28 ( .A(n108), .B(n106), .CO(n38), .S(n39) );
  CMPR42X1 U29 ( .A(n109), .B(n107), .C(a[5]), .D(a[7]), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U30 ( .A(a[4]), .B(a[6]), .CI(n46), .CO(n43), .S(n44) );
  ADDFXL U33 ( .A(a[3]), .B(n109), .CI(a[5]), .CO(n47), .S(n48) );
  BUFX6 U51 ( .A(a[1]), .Y(n99) );
  CLKBUFX3 U52 ( .A(a[2]), .Y(n100) );
  CLKBUFX2 U53 ( .A(n99), .Y(product[1]) );
  INVXL U54 ( .A(n99), .Y(n109) );
  CLKBUFX3 U55 ( .A(a[0]), .Y(product[0]) );
  CLKINVX1 U56 ( .A(a[4]), .Y(n106) );
  CLKINVX1 U57 ( .A(n100), .Y(n108) );
  CLKINVX1 U58 ( .A(a[3]), .Y(n107) );
  CLKINVX1 U59 ( .A(a[6]), .Y(n104) );
  CLKINVX1 U60 ( .A(a[5]), .Y(n105) );
  CLKINVX1 U61 ( .A(a[7]), .Y(n103) );
  XOR2X1 U62 ( .A(n104), .B(n110), .Y(product[16]) );
  XOR2X1 U63 ( .A(n2), .B(a[7]), .Y(n110) );
  XOR2X1 U64 ( .A(a[4]), .B(a[0]), .Y(n50) );
  NAND2X1 U65 ( .A(a[0]), .B(n106), .Y(n49) );
  XOR2X1 U66 ( .A(n108), .B(a[0]), .Y(n46) );
  NAND2X1 U67 ( .A(a[0]), .B(n100), .Y(n45) );
endmodule


module imgproc_DW_mult_uns_9 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[3]), .Y(n74) );
  CLKINVX1 U37 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U38 ( .A(a[1]), .Y(n76) );
  CLKBUFX3 U39 ( .A(a[0]), .Y(product_3_) );
  CLKINVX1 U40 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U41 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U42 ( .A(a[6]), .Y(n71) );
  CLKINVX1 U43 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U44 ( .A(a[7]), .Y(n70) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW_mult_uns_7 ( a, product );
  input [7:0] a;
  output [19:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n89, n90,
         n91, n92, n93, n94, n95, n96, n97;

  ADDFXL U3 ( .A(n90), .B(a[5]), .CI(n3), .CO(n2), .S(product[18]) );
  ADDFXL U4 ( .A(n20), .B(n91), .CI(n4), .CO(n3), .S(product[17]) );
  ADDFXL U5 ( .A(n21), .B(n22), .CI(n5), .CO(n4), .S(product[16]) );
  ADDFXL U6 ( .A(n23), .B(n24), .CI(n6), .CO(n5), .S(product[15]) );
  ADDFXL U7 ( .A(n26), .B(n25), .CI(n7), .CO(n6), .S(product[14]) );
  ADDFXL U8 ( .A(n27), .B(n28), .CI(n8), .CO(n7), .S(product[13]) );
  ADDFXL U9 ( .A(n29), .B(n30), .CI(n9), .CO(n8), .S(product[12]) );
  ADDFXL U10 ( .A(n31), .B(n32), .CI(n10), .CO(n9), .S(product[11]) );
  ADDFXL U11 ( .A(n33), .B(a[4]), .CI(n11), .CO(n10), .S(product[10]) );
  ADDFXL U12 ( .A(a[3]), .B(a[0]), .CI(n12), .CO(n11), .S(product[9]) );
  ADDHXL U13 ( .A(a[2]), .B(n13), .CO(n12), .S(product[8]) );
  ADDFXL U14 ( .A(a[7]), .B(a[1]), .CI(n14), .CO(n13), .S(product[7]) );
  ADDHXL U15 ( .A(a[0]), .B(a[6]), .CO(n14), .S(product[6]) );
  ADDHXL U19 ( .A(n89), .B(a[4]), .CO(n20), .S(n21) );
  ADDHXL U20 ( .A(n90), .B(a[3]), .CO(n22), .S(n23) );
  ADDHXL U21 ( .A(n91), .B(a[2]), .CO(n24), .S(n25) );
  ADDFXL U22 ( .A(a[1]), .B(n92), .CI(a[7]), .CO(n26), .S(n27) );
  ADDFXL U23 ( .A(a[0]), .B(n93), .CI(a[6]), .CO(n28), .S(n29) );
  ADDHXL U24 ( .A(n94), .B(a[5]), .CO(n30), .S(n31) );
  ADDHXL U25 ( .A(n96), .B(n95), .CO(n32), .S(n33) );
  CLKBUFX3 U41 ( .A(a[1]), .Y(product[1]) );
  CLKBUFX3 U42 ( .A(a[2]), .Y(product[2]) );
  CLKBUFX3 U43 ( .A(a[3]), .Y(product[3]) );
  CLKBUFX3 U44 ( .A(a[0]), .Y(product[0]) );
  CLKBUFX3 U45 ( .A(a[4]), .Y(product[4]) );
  CLKBUFX3 U46 ( .A(a[5]), .Y(product[5]) );
  CLKINVX1 U47 ( .A(a[1]), .Y(n95) );
  CLKINVX1 U48 ( .A(a[0]), .Y(n96) );
  CLKINVX1 U49 ( .A(a[2]), .Y(n94) );
  CLKINVX1 U50 ( .A(a[3]), .Y(n93) );
  CLKINVX1 U51 ( .A(a[4]), .Y(n92) );
  CLKINVX1 U52 ( .A(a[6]), .Y(n90) );
  CLKINVX1 U53 ( .A(a[5]), .Y(n91) );
  CLKINVX1 U54 ( .A(a[7]), .Y(n89) );
  XOR2X1 U55 ( .A(n90), .B(n97), .Y(product[19]) );
  XOR2X1 U56 ( .A(n2), .B(a[7]), .Y(n97) );
endmodule


module imgproc_DW_mult_uns_5 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U37 ( .A(a[1]), .Y(n76) );
  CLKBUFX3 U38 ( .A(a[0]), .Y(product_3_) );
  CLKINVX1 U39 ( .A(a[3]), .Y(n74) );
  CLKINVX1 U40 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U41 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U42 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U43 ( .A(a[6]), .Y(n71) );
  CLKINVX1 U44 ( .A(a[7]), .Y(n70) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW_mult_uns_3 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U37 ( .A(a[1]), .Y(n76) );
  CLKINVX1 U38 ( .A(a[3]), .Y(n74) );
  CLKBUFX3 U39 ( .A(a[0]), .Y(product_3_) );
  CLKINVX1 U40 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U41 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U42 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U43 ( .A(a[6]), .Y(n71) );
  CLKINVX1 U44 ( .A(a[7]), .Y(n70) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW_mult_uns_2 ( a, product );
  input [7:0] a;
  output [16:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n101, n102, n103, n104, n105, n106, n107, n108;

  ADDFXL U3 ( .A(n19), .B(n102), .CI(n3), .CO(n2), .S(product[15]) );
  ADDFXL U4 ( .A(n21), .B(n20), .CI(n4), .CO(n3), .S(product[14]) );
  ADDFXL U5 ( .A(n23), .B(n22), .CI(n5), .CO(n4), .S(product[13]) );
  ADDFXL U6 ( .A(n25), .B(n24), .CI(n6), .CO(n5), .S(product[12]) );
  ADDFXL U7 ( .A(n26), .B(n29), .CI(n7), .CO(n6), .S(product[11]) );
  ADDFXL U8 ( .A(n30), .B(n34), .CI(n8), .CO(n7), .S(product[10]) );
  ADDFXL U9 ( .A(n36), .B(n35), .CI(n9), .CO(n8), .S(product[9]) );
  ADDFXL U10 ( .A(n37), .B(n41), .CI(n10), .CO(n9), .S(product[8]) );
  ADDFXL U11 ( .A(n43), .B(n42), .CI(n11), .CO(n10), .S(product[7]) );
  ADDFXL U12 ( .A(n44), .B(n47), .CI(n12), .CO(n11), .S(product[6]) );
  ADDFXL U13 ( .A(n48), .B(n49), .CI(n13), .CO(n12), .S(product[5]) );
  ADDFXL U14 ( .A(n50), .B(a[2]), .CI(n14), .CO(n13), .S(product[4]) );
  ADDFXL U15 ( .A(a[3]), .B(a[1]), .CI(n15), .CO(n14), .S(product[3]) );
  ADDHXL U19 ( .A(n101), .B(a[5]), .CO(n19), .S(n20) );
  ADDFXL U20 ( .A(n102), .B(a[7]), .CI(a[4]), .CO(n21), .S(n22) );
  ADDFXL U21 ( .A(a[3]), .B(a[6]), .CI(n27), .CO(n23), .S(n24) );
  ADDFXL U22 ( .A(n31), .B(a[2]), .CI(n28), .CO(n25), .S(n26) );
  ADDHXL U23 ( .A(n101), .B(n103), .CO(n27), .S(n28) );
  ADDFXL U24 ( .A(n33), .B(a[1]), .CI(n32), .CO(n29), .S(n30) );
  ADDHXL U25 ( .A(n102), .B(n104), .CO(n31), .S(n32) );
  CMPR42X1 U26 ( .A(n105), .B(n103), .C(a[0]), .D(a[7]), .ICI(n38), .S(n35), 
        .ICO(n33), .CO(n34) );
  ADDFXL U27 ( .A(n40), .B(a[6]), .CI(n39), .CO(n36), .S(n37) );
  ADDHXL U28 ( .A(n106), .B(n104), .CO(n38), .S(n39) );
  CMPR42X1 U29 ( .A(n107), .B(n105), .C(a[5]), .D(a[7]), .ICI(n45), .S(n42), 
        .ICO(n40), .CO(n41) );
  ADDFXL U30 ( .A(a[4]), .B(a[6]), .CI(n46), .CO(n43), .S(n44) );
  ADDFXL U33 ( .A(a[3]), .B(n107), .CI(a[5]), .CO(n47), .S(n48) );
  ADDHX1 U51 ( .A(a[0]), .B(a[2]), .CO(n15), .S(product[2]) );
  CLKBUFX2 U52 ( .A(a[1]), .Y(product[1]) );
  INVXL U53 ( .A(a[1]), .Y(n107) );
  XOR2XL U54 ( .A(a[4]), .B(a[0]), .Y(n50) );
  NAND2XL U55 ( .A(a[0]), .B(n104), .Y(n49) );
  INVXL U56 ( .A(a[2]), .Y(n106) );
  XOR2XL U57 ( .A(n106), .B(a[0]), .Y(n46) );
  NAND2XL U58 ( .A(a[0]), .B(a[2]), .Y(n45) );
  CLKBUFX3 U59 ( .A(a[0]), .Y(product[0]) );
  CLKINVX1 U60 ( .A(a[4]), .Y(n104) );
  CLKINVX1 U61 ( .A(a[3]), .Y(n105) );
  CLKINVX1 U62 ( .A(a[6]), .Y(n102) );
  CLKINVX1 U63 ( .A(a[5]), .Y(n103) );
  CLKINVX1 U64 ( .A(a[7]), .Y(n101) );
  XOR2X1 U65 ( .A(n102), .B(n108), .Y(product[16]) );
  XOR2X1 U66 ( .A(n2), .B(a[7]), .Y(n108) );
endmodule


module imgproc_DW_mult_uns_1 ( a, product_15_, product_14_, product_13_, 
        product_12_, product_11_, product_10_, product_9_, product_8_, 
        product_7_, product_6_, product_5_, product_4_, product_3_ );
  input [7:0] a;
  output product_15_, product_14_, product_13_, product_12_, product_11_,
         product_10_, product_9_, product_8_, product_7_, product_6_,
         product_5_, product_4_, product_3_;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n70, n71, n72, n73, n74,
         n75, n76, n77, n78;

  ADDFXL U4 ( .A(n13), .B(a[5]), .CI(n3), .CO(n2), .S(product_13_) );
  ADDFXL U5 ( .A(n14), .B(n15), .CI(n4), .CO(n3), .S(product_12_) );
  ADDFXL U6 ( .A(n17), .B(n16), .CI(n5), .CO(n4), .S(product_11_) );
  ADDFXL U7 ( .A(n18), .B(n19), .CI(n6), .CO(n5), .S(product_10_) );
  ADDFXL U8 ( .A(n20), .B(n21), .CI(n7), .CO(n6), .S(product_9_) );
  ADDFXL U9 ( .A(n22), .B(n23), .CI(n8), .CO(n7), .S(product_8_) );
  ADDFXL U10 ( .A(n24), .B(n25), .CI(n9), .CO(n8), .S(product_7_) );
  ADDFXL U11 ( .A(n26), .B(n75), .CI(n10), .CO(n9), .S(product_6_) );
  ADDFXL U12 ( .A(n77), .B(a[2]), .CI(n11), .CO(n10), .S(product_5_) );
  ADDHXL U13 ( .A(n76), .B(n77), .CO(n11), .S(product_4_) );
  ADDFXL U19 ( .A(n72), .B(n70), .CI(a[2]), .CO(n17), .S(n18) );
  ADDFXL U20 ( .A(n73), .B(n71), .CI(a[1]), .CO(n19), .S(n20) );
  ADDFXL U21 ( .A(n74), .B(n72), .CI(a[0]), .CO(n21), .S(n22) );
  ADDHXL U22 ( .A(n73), .B(n75), .CO(n23), .S(n24) );
  ADDHXL U23 ( .A(n74), .B(n76), .CO(n25), .S(n26) );
  CLKINVX1 U36 ( .A(a[0]), .Y(n77) );
  CLKINVX1 U37 ( .A(a[1]), .Y(n76) );
  CLKBUFX3 U38 ( .A(a[0]), .Y(product_3_) );
  CLKINVX1 U39 ( .A(a[3]), .Y(n74) );
  CLKINVX1 U40 ( .A(a[2]), .Y(n75) );
  CLKINVX1 U41 ( .A(a[4]), .Y(n73) );
  CLKINVX1 U42 ( .A(a[5]), .Y(n72) );
  CLKINVX1 U43 ( .A(a[6]), .Y(n71) );
  CLKINVX1 U44 ( .A(a[7]), .Y(n70) );
  XNOR2X1 U45 ( .A(n70), .B(n78), .Y(product_15_) );
  NOR2X1 U46 ( .A(a[6]), .B(n2), .Y(n78) );
  XNOR2X1 U47 ( .A(n2), .B(a[6]), .Y(product_14_) );
  XNOR2X1 U48 ( .A(n71), .B(a[3]), .Y(n16) );
  NAND2X1 U49 ( .A(a[6]), .B(n74), .Y(n15) );
  XNOR2X1 U50 ( .A(n70), .B(a[4]), .Y(n14) );
  NAND2X1 U51 ( .A(a[7]), .B(n73), .Y(n13) );
endmodule


module imgproc_DW01_add_19 ( A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, 
        A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_16_, 
        B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, 
        B_4_, B_3_, B_2_, B_1_, B_0_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, 
        SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_,
         A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_16_, B_15_, B_14_, B_13_,
         B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_,
         B_1_, B_0_;
  output SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_,
         SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_,
         SUM_2_, SUM_1_, SUM_0_;
  wire   n1;
  wire   [16:2] carry;

  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(SUM_17_), .S(
        SUM_16_) );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_16 ( A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, 
        A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, 
        A_0_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, 
        B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_19_, 
        SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, 
        SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, 
        SUM_2_, SUM_1_, SUM_0_ );
  input A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_,
         A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_18_, B_17_,
         B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_,
         B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_,
         SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_,
         SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   n1;
  wire   [18:2] carry;

  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(SUM_19_), .S(
        SUM_18_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_15 ( A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, 
        A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, 
        A_1_, A_0_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, 
        B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, 
        B_0_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, 
        SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_,
         A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_,
         SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_,
         SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   n1;
  wire   [19:2] carry;

  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(SUM_20_), .S(
        SUM_19_) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_14 ( A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, 
        A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, 
        A_1_, A_0_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, 
        B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, 
        B_0_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, 
        SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_,
         A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_,
         SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_,
         SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   n1;
  wire   [19:2] carry;

  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry[19]), .CO(SUM_20_), .S(
        SUM_19_) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_13 ( A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, 
        A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, 
        A_2_, A_1_, A_0_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, 
        B_2_, B_1_, B_0_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_,
         A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_,
         B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_,
         B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   carry_20_, carry_19_, carry_18_, carry_17_, carry_16_, carry_15_,
         carry_14_, carry_13_, carry_12_, carry_11_, carry_10_, carry_9_,
         carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_,
         n1;

  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(SUM_21_), .S(
        SUM_20_) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry_5_), .CO(carry_6_), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry_4_), .CO(carry_5_), .S(SUM_4_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry_2_), .CO(carry_3_), .S(SUM_2_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry_3_), .CO(carry_4_), .S(SUM_3_)
         );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry_2_), .S(SUM_1_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry_6_), .CO(carry_7_), .S(SUM_6_)
         );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_9 ( A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, 
        A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, 
        A_0_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, 
        B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_19_, 
        SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, 
        SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, 
        SUM_2_, SUM_1_, SUM_0_ );
  input A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_,
         A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_18_, B_17_,
         B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_,
         B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_,
         SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_,
         SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   carry_18_, carry_17_, carry_16_, carry_15_, carry_14_, carry_13_,
         carry_12_, carry_11_, carry_10_, carry_9_, carry_8_, carry_7_,
         carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1;

  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(SUM_19_), .S(
        SUM_18_) );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry_2_), .S(SUM_1_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry_2_), .CO(carry_3_), .S(SUM_2_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry_3_), .CO(carry_4_), .S(SUM_3_)
         );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry_5_), .CO(carry_6_), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry_4_), .CO(carry_5_), .S(SUM_4_)
         );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry_6_), .CO(carry_7_), .S(SUM_6_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_8 ( A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, 
        A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, 
        A_0_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, 
        B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_, SUM_19_, 
        SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, 
        SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, 
        SUM_2_, SUM_1_, SUM_0_ );
  input A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_,
         A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_18_, B_17_,
         B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_,
         B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, SUM_13_,
         SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, SUM_5_,
         SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   n1;
  wire   [18:2] carry;

  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry[18]), .CO(SUM_19_), .S(
        SUM_18_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry[2]), .S(SUM_1_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry[13]), .CO(carry[14]), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry[12]), .CO(carry[13]), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry[11]), .CO(carry[12]), .S(
        SUM_11_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry[10]), .CO(carry[11]), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry[9]), .CO(carry[10]), .S(SUM_9_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry[8]), .CO(carry[9]), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry[7]), .CO(carry[8]), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry[6]), .CO(carry[7]), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry[5]), .CO(carry[6]), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry[4]), .CO(carry[5]), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry[3]), .CO(carry[4]), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry[2]), .CO(carry[3]), .S(SUM_2_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_7 ( A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, 
        A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, 
        A_1_, A_0_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, 
        B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, 
        B_0_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_, 
        SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_, 
        SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_, A_10_,
         A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_, B_19_,
         B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_, B_9_,
         B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_, SUM_14_,
         SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_, SUM_6_,
         SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   carry_19_, carry_18_, carry_17_, carry_16_, carry_15_, carry_14_,
         carry_13_, carry_12_, carry_11_, carry_10_, carry_9_, carry_8_,
         carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_, n1;

  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(SUM_20_), .S(
        SUM_19_) );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry_2_), .S(SUM_1_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry_6_), .CO(carry_7_), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry_5_), .CO(carry_6_), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry_4_), .CO(carry_5_), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry_3_), .CO(carry_4_), .S(SUM_3_)
         );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry_2_), .CO(carry_3_), .S(SUM_2_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_4 ( A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, 
        A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, 
        A_2_, A_1_, A_0_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, 
        B_2_, B_1_, B_0_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, 
        SUM_15_, SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, 
        SUM_7_, SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_ );
  input A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_, A_11_,
         A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_, A_0_,
         B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_,
         B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  output SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_, SUM_15_,
         SUM_14_, SUM_13_, SUM_12_, SUM_11_, SUM_10_, SUM_9_, SUM_8_, SUM_7_,
         SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_, SUM_0_;
  wire   carry_20_, carry_19_, carry_18_, carry_17_, carry_16_, carry_15_,
         carry_14_, carry_13_, carry_12_, carry_11_, carry_10_, carry_9_,
         carry_8_, carry_7_, carry_6_, carry_5_, carry_4_, carry_3_, carry_2_,
         n1;

  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM_19_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM_18_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM_16_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(SUM_21_), .S(
        SUM_20_) );
  ADDFXL U1_1 ( .A(A_1_), .B(B_1_), .CI(n1), .CO(carry_2_), .S(SUM_1_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM_17_) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM_15_) );
  ADDFXL U1_2 ( .A(A_2_), .B(B_2_), .CI(carry_2_), .CO(carry_3_), .S(SUM_2_)
         );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM_14_) );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM_13_) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM_12_) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM_11_) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM_10_) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM_9_)
         );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM_8_)
         );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM_7_)
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry_6_), .CO(carry_7_), .S(SUM_6_)
         );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry_5_), .CO(carry_6_), .S(SUM_5_)
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(carry_4_), .CO(carry_5_), .S(SUM_4_)
         );
  ADDFXL U1_3 ( .A(A_3_), .B(B_3_), .CI(carry_3_), .CO(carry_4_), .S(SUM_3_)
         );
  AND2X2 U1 ( .A(B_0_), .B(A_0_), .Y(n1) );
  XOR2X1 U2 ( .A(B_0_), .B(A_0_), .Y(SUM_0_) );
endmodule


module imgproc_DW01_add_3 ( SUM, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, 
        A_15_, A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, 
        A_4_, A_3_, B_21_, B_20_, B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, 
        B_2_, B_1_, B_0_ );
  output [22:0] SUM;
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, B_21_, B_20_,
         B_19_, B_18_, B_17_, B_16_, B_15_, B_14_, B_13_, B_12_, B_11_, B_10_,
         B_9_, B_8_, B_7_, B_6_, B_5_, B_4_, B_3_, B_2_, B_1_, B_0_;
  wire   carry_21_, carry_20_, carry_19_, carry_18_, carry_17_, carry_16_,
         carry_15_, carry_14_, carry_13_, carry_12_, carry_11_, carry_10_,
         carry_9_, carry_8_, carry_7_, carry_6_, carry_5_, n1;

  ADDFXL U1_20 ( .A(A_20_), .B(B_20_), .CI(carry_20_), .CO(carry_21_), .S(
        SUM[20]) );
  ADDFXL U1_21 ( .A(A_21_), .B(B_21_), .CI(carry_21_), .CO(SUM[22]), .S(
        SUM[21]) );
  ADDFXL U1_5 ( .A(A_5_), .B(B_5_), .CI(carry_5_), .CO(carry_6_), .S(SUM[5])
         );
  ADDFXL U1_4 ( .A(A_4_), .B(B_4_), .CI(n1), .CO(carry_5_), .S(SUM[4]) );
  ADDFXL U1_18 ( .A(A_18_), .B(B_18_), .CI(carry_18_), .CO(carry_19_), .S(
        SUM[18]) );
  ADDFXL U1_8 ( .A(A_8_), .B(B_8_), .CI(carry_8_), .CO(carry_9_), .S(SUM[8])
         );
  ADDFXL U1_19 ( .A(A_19_), .B(B_19_), .CI(carry_19_), .CO(carry_20_), .S(
        SUM[19]) );
  ADDFXL U1_7 ( .A(A_7_), .B(B_7_), .CI(carry_7_), .CO(carry_8_), .S(SUM[7])
         );
  ADDFXL U1_6 ( .A(A_6_), .B(B_6_), .CI(carry_6_), .CO(carry_7_), .S(SUM[6])
         );
  ADDFXL U1_13 ( .A(A_13_), .B(B_13_), .CI(carry_13_), .CO(carry_14_), .S(
        SUM[13]) );
  ADDFXL U1_17 ( .A(A_17_), .B(B_17_), .CI(carry_17_), .CO(carry_18_), .S(
        SUM[17]) );
  ADDFXL U1_16 ( .A(A_16_), .B(B_16_), .CI(carry_16_), .CO(carry_17_), .S(
        SUM[16]) );
  ADDFXL U1_15 ( .A(A_15_), .B(B_15_), .CI(carry_15_), .CO(carry_16_), .S(
        SUM[15]) );
  ADDFXL U1_14 ( .A(A_14_), .B(B_14_), .CI(carry_14_), .CO(carry_15_), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A_12_), .B(B_12_), .CI(carry_12_), .CO(carry_13_), .S(
        SUM[12]) );
  ADDFXL U1_11 ( .A(A_11_), .B(B_11_), .CI(carry_11_), .CO(carry_12_), .S(
        SUM[11]) );
  ADDFXL U1_10 ( .A(A_10_), .B(B_10_), .CI(carry_10_), .CO(carry_11_), .S(
        SUM[10]) );
  ADDFXL U1_9 ( .A(A_9_), .B(B_9_), .CI(carry_9_), .CO(carry_10_), .S(SUM[9])
         );
  AND2X2 U1 ( .A(B_3_), .B(A_3_), .Y(n1) );
  CLKBUFX3 U2 ( .A(B_2_), .Y(SUM[2]) );
  CLKBUFX3 U3 ( .A(B_0_), .Y(SUM[0]) );
  CLKBUFX3 U4 ( .A(B_1_), .Y(SUM[1]) );
  XOR2X1 U5 ( .A(B_3_), .B(A_3_), .Y(SUM[3]) );
endmodule


module imgproc_DW01_add_2 ( B, A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, 
        A_14_, A_13_, A_12_, A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, 
        A_3_, A_2_, A_1_, A_0_, SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, 
        SUM_17_, SUM_16_, SUM_15_, SUM_14_ );
  input [22:0] B;
  input A_21_, A_20_, A_19_, A_18_, A_17_, A_16_, A_15_, A_14_, A_13_, A_12_,
         A_11_, A_10_, A_9_, A_8_, A_7_, A_6_, A_5_, A_4_, A_3_, A_2_, A_1_,
         A_0_;
  output SUM_22_, SUM_21_, SUM_20_, SUM_19_, SUM_18_, SUM_17_, SUM_16_,
         SUM_15_, SUM_14_;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [22:14] carry;

  ADDFXL U1_15 ( .A(A_15_), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM_15_) );
  ADDFXL U1_19 ( .A(A_19_), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM_19_) );
  ADDFXL U1_17 ( .A(A_17_), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM_17_) );
  ADDFXL U1_21 ( .A(A_21_), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM_21_) );
  ADDFXL U1_18 ( .A(A_18_), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM_18_) );
  ADDFXL U1_16 ( .A(A_16_), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM_16_) );
  ADDFXL U1_14 ( .A(A_14_), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM_14_) );
  ADDFXL U1_20 ( .A(A_20_), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM_20_) );
  OAI21XL U1 ( .A0(A_13_), .A1(n1), .B0(B[13]), .Y(n2) );
  XOR2X1 U2 ( .A(B[22]), .B(carry[22]), .Y(SUM_22_) );
  OAI2BB1X1 U3 ( .A0N(n1), .A1N(A_13_), .B0(n2), .Y(carry[14]) );
  OAI2BB1X1 U4 ( .A0N(n3), .A1N(A_12_), .B0(n4), .Y(n1) );
  OAI21XL U5 ( .A0(A_12_), .A1(n3), .B0(B[12]), .Y(n4) );
  OAI2BB1X1 U6 ( .A0N(n5), .A1N(A_11_), .B0(n6), .Y(n3) );
  OAI21XL U7 ( .A0(A_11_), .A1(n5), .B0(B[11]), .Y(n6) );
  OAI2BB1X1 U8 ( .A0N(n7), .A1N(A_10_), .B0(n8), .Y(n5) );
  OAI21XL U9 ( .A0(A_10_), .A1(n7), .B0(B[10]), .Y(n8) );
  OAI2BB1X1 U10 ( .A0N(n9), .A1N(A_9_), .B0(n10), .Y(n7) );
  OAI21XL U11 ( .A0(A_9_), .A1(n9), .B0(B[9]), .Y(n10) );
  OAI2BB1X1 U12 ( .A0N(n11), .A1N(A_8_), .B0(n12), .Y(n9) );
  OAI21XL U13 ( .A0(A_8_), .A1(n11), .B0(B[8]), .Y(n12) );
  OAI2BB1X1 U14 ( .A0N(n13), .A1N(A_7_), .B0(n14), .Y(n11) );
  OAI21XL U15 ( .A0(A_7_), .A1(n13), .B0(B[7]), .Y(n14) );
  OAI2BB1X1 U16 ( .A0N(n15), .A1N(A_6_), .B0(n16), .Y(n13) );
  OAI21XL U17 ( .A0(A_6_), .A1(n15), .B0(B[6]), .Y(n16) );
  OAI2BB1X1 U18 ( .A0N(n17), .A1N(A_5_), .B0(n18), .Y(n15) );
  OAI21XL U19 ( .A0(A_5_), .A1(n17), .B0(B[5]), .Y(n18) );
  OAI2BB1X1 U20 ( .A0N(n19), .A1N(A_4_), .B0(n20), .Y(n17) );
  OAI21XL U21 ( .A0(A_4_), .A1(n19), .B0(B[4]), .Y(n20) );
  OAI2BB1X1 U22 ( .A0N(n21), .A1N(A_3_), .B0(n22), .Y(n19) );
  OAI21XL U23 ( .A0(A_3_), .A1(n21), .B0(B[3]), .Y(n22) );
  OAI2BB1X1 U24 ( .A0N(n23), .A1N(A_2_), .B0(n24), .Y(n21) );
  OAI21XL U25 ( .A0(A_2_), .A1(n23), .B0(B[2]), .Y(n24) );
  OAI2BB1X1 U26 ( .A0N(A_1_), .A1N(B[1]), .B0(n25), .Y(n23) );
  OAI211X1 U27 ( .A0(A_1_), .A1(B[1]), .B0(A_0_), .C0(B[0]), .Y(n25) );
endmodule


module imgproc_DW01_inc_5 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  XOR2X1 U1 ( .A(carry[7]), .B(A[7]), .Y(SUM[7]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module imgproc ( clk, rst, orig_data, orig_ready, request, orig_addr, 
        imgproc_ready, imgproc_addr, imgproc_data, finish );
  input [7:0] orig_data;
  output [13:0] orig_addr;
  output [13:0] imgproc_addr;
  output [7:0] imgproc_data;
  input clk, rst, orig_ready;
  output request, imgproc_ready, finish;
  wire   n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         next_imgproc_ready, next_finish, next_request, N114, N115, N116, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1270, N1271, N1272, N1273, N1274, N1275,
         N1276, N1277, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289,
         N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245, N2246, N2250,
         N2251, N2252, N2253, N2254, N2255, N2256, N2257, N2274, N2275, N2276,
         N2277, N2278, N2279, N2280, N2281, N2282, N2283, N2284, N2285, N2286,
         N2287, n1640, n1650, n1660, n1680, n1690, n1700, n1710, n1720, n1730,
         n1740, n1750, n1760, n1770, n1780, n1790, n1800, n1810, n1820, n1830,
         n1840, n1850, n1860, n1870, n1880, n1890, n1900, n1910, n1920, n1930,
         n1940, n1950, n1960, n1970, n1980, n1990, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n224, n225, n226, n227, n228, n229, n230, n231, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n304,
         n305, n306, n307, n308, n309, n310, n311, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n6680,
         n6690, n6700, n6710, n6720, n6730, n6740, n6750, n6760, n6770, n6780,
         n6790, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, N2237, N2236, N2235, N2234, N2233, N2232, N2231,
         N2230, N2229, N2228, N2227, N2226, N2221, N2220, N2219, N2218, N2217,
         N2216, N2215, N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207,
         N2206, N2205, N2204, N2203, N2202, N2201, N2200, N2199, N2198, N2197,
         N2196, N2195, N2194, N2193, N2192, N2191, N2190, N2189, N2185, N2184,
         N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174,
         N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164,
         N2163, N2162, N2161, N2160, N2159, N2158, N2157, N2156, N2155, N2154,
         N2153, N2152, N2151, N2150, N2149, N2148, N2147, N2146, N2140, N2139,
         N2138, N2137, N2136, N2135, N2134, N2133, N2132, N2131, N2130, N2129,
         N2128, N2127, N2126, N2122, N2121, N2120, N2119, N2118, N2117, N2116,
         N2115, N2114, N2113, N2112, N2111, N2110, N2104, N2103, N2102, N2101,
         N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, N2092, N2091,
         N2090, N2089, N2088, N2087, N2086, N2085, N2084, N2083, N2082, N2081,
         N2080, N2079, N2078, N2077, N2076, N2075, N2074, N2073, N2072, N2067,
         N2066, N2065, N2064, N2063, N2062, N2061, N2060, N2059, N2058, N2057,
         N2056, N2055, N2054, N2053, N2052, N2051, N2050, N2049, N2048, N2047,
         N2046, N2045, N2044, N2043, N2042, N2041, N2040, N2039, N2038, N2037,
         N2036, N2035, N2030, N2029, N2028, N2027, N2026, N2025, N2024, N2023,
         N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014, N2013,
         N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004, N2003,
         N2002, N2001, N2000, N1999, N1998, N1997, N1996, N1995, N1994, N1993,
         N1992, N1991, N19900, N1983, N1982, N1981, N19800, N1979, N1978,
         N1977, N1976, N1975, N1974, N1973, N1972, N1971, N19700, N1966, N1965,
         N1964, N1963, N1962, N1961, N19600, N1959, N1958, N1957, N1956, N1955,
         N1954, N1953, N1952, N1951, N19500, N1949, N1948, N1947, N19400,
         N1939, N1938, N1937, N1936, N1935, N1934, N1933, N1932, N1931, N19300,
         N1929, N1928, N1927, N1923, N1922, N1921, N19200, N1919, N1918, N1917,
         N1916, N1915, N1914, N1913, N1912, N1911, N19100, N1909, N1908, N1907,
         N1906, N1905, N1901, N19000, N1899, N1898, N1897, N1896, N1895, N1894,
         N1893, N1892, N1891, N18900, N1889, N1888, N1887, N1886, N1885, N1884,
         N1883, N1882, N1881, N18800, N1879, N1878, N1877, N1876, N1875, N1874,
         N1873, N1872, N1871, N18700, N1869, N1863, N1862, N1861, N18600,
         N1859, N1858, N1857, N1856, N1855, N1854, N1853, N1852, N1851, N18500,
         N1849, N1848, N1847, N1846, N1845, N1844, N1843, N1842, N1841, N18400,
         N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, N18300,
         N1829, N1828, N1827, N1826, N18200, N1819, N1818, N1817, N1816, N1815,
         N1814, N1813, N1812, N1811, N18100, N1809, N1808, N1807, N1806, N1805,
         N1804, N1803, N1802, N1801, N18000, N1799, N1798, N1797, N1796, N1795,
         N1794, N1793, N1792, N1791, N17900, N1789, N1788, N1787, N1786, N1785,
         N1784, N1783, N17800, N1779, N1778, N1777, N1776, N1775, N1774, N1773,
         N1772, N1771, N17700, N1769, N1768, N1767, N1766, N1765, N1764, N1763,
         N1759, N1758, N1757, N1756, N1755, N1754, N1753, N1752, N1751, N17500,
         N1749, N1748, N1747, N1746, N1745, N1744, N1743, N1742, N1736, N1735,
         N1734, N1733, N1732, N1731, N17300, N1729, N1728, N1727, N1726, N1725,
         N1724, N1723, N1722, N1721, N17200, N1719, N1718, N1717, N1716, N1715,
         N1714, N1713, N1712, N1711, N17100, N1709, N1708, N1707, N1706, N1705,
         N1704, N1703, N1702, N1701, N17000, N1699, N1698, N1697, N1696, N1694,
         N1693, N1692, N1691, N16900, N1689, N1688, N1687, N1686, N1685, N1684,
         N1683, N1682, N1681, N16800, N1679, N1678, N1677, N1676, N1675, N1674,
         N1673, N1672, N1671, N1670, N1669, N1668, N1667, N1666, N1665, N1664,
         N1663, N1662, N1661, N16600, N1659, N1658, N1657, N1656, N1646, N1645,
         N1644, N1643, N1642, N1641, N16400, N1639, N1638, N1637, N1636, N1635,
         N1634, N1632, N1631, N1630, N1629, N1628, N1627, N1626, N1625, N1624,
         N1623, N1622, N1621, N1620, N1607, N1606, N1605, N1604, N1603, N1602,
         N1601, N1600, N1599, N1598, N1597, N1596, N1595, N1593, N1592, N1591,
         N1590, N1589, N1588, N1587, N1586, N1585, N1584, N1583, N1582, N1581,
         N1580, N1579, N1578, N1577, N1576, N1575, N1568, N1567, N1566, N1565,
         N1564, N1563, N1562, N1561, N1560, N1559, N1558, N1557, N1556, N1555,
         N1551, N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542,
         N1541, N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532,
         N1526, N1525, N1524, N1523, N1522, N1521, N1520, N1519, N1518, N1517,
         N1516, N1515, N1514, N1513, N1509, N1508, N1507, N1506, N1505, N1504,
         N1503, N1502, N1501, N1500, N1499, N1498, N1497, N1496, N1495, N1494,
         N1493, N1492, N1491, N1487, N1486, N1485, N1484, N1483, N1482, N1481,
         N1480, N1479, N1478, N1477, N1476, N1475, N1474, N1473, N1472, N1471,
         N1470, N1469, N1468, N1467, N1466, N1465, N1464, N1463, N1462, N1461,
         N1460, N1459, N1458, N1457, N1433, N1432, N1431, N1430, N1429, N1428,
         N1427, N1426, N1425, N1424, N1423, N1422, N1401, N1400, N1399, N1398,
         N1397, N1396, N1395, N1394, N1393, N1392, N1391, N1390, N1389, N1367,
         N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357,
         N1356, N1355, N1354, N1353, N1352, N1351, N1333, N1332, N1331, N1330,
         N1329, N1328, N1327, N1326, N1325, N1324, N1323, N1322, N1321, N13170,
         N13160, N13150, N13140, N13130, N13120, N13110, N13100, N13090,
         N13080, N13070, N13060, sub_203_carry_2_, sub_203_carry_3_,
         sub_203_carry_4_, sub_203_carry_5_, sub_203_carry_6_,
         sub_203_carry_7_, sub_203_carry_8_, sub_203_carry_10_,
         sub_203_carry_11_, sub_203_carry_12_, sub_203_carry_13_,
         sub_139_carry_3_, sub_139_carry_8_, sub_139_carry_9_,
         sub_139_carry_11_, sub_139_carry_12_, sub_139_carry_13_,
         r652_carry_8_, r652_carry_9_, r652_carry_11_, r652_carry_12_,
         r652_carry_13_, add_9_root_add_0_root_add_245_5_carry_3_,
         add_9_root_add_0_root_add_245_5_carry_4_,
         add_9_root_add_0_root_add_245_5_carry_5_,
         add_9_root_add_0_root_add_245_5_carry_6_,
         add_9_root_add_0_root_add_245_5_carry_7_,
         add_9_root_add_0_root_add_245_5_carry_8_,
         add_9_root_add_0_root_add_245_5_carry_9_,
         add_9_root_add_0_root_add_245_5_carry_10_,
         add_9_root_add_0_root_add_245_5_carry_11_,
         add_9_root_add_0_root_add_245_5_carry_12_,
         add_9_root_add_0_root_add_245_5_carry_13_,
         add_9_root_add_0_root_add_245_5_carry_14_,
         add_9_root_add_0_root_add_245_5_carry_15_,
         add_9_root_add_0_root_add_245_5_B_1_,
         add_9_root_add_0_root_add_245_5_B_2_,
         add_9_root_add_0_root_add_245_5_B_3_,
         add_9_root_add_0_root_add_245_5_B_4_,
         add_9_root_add_0_root_add_245_5_B_5_,
         add_9_root_add_0_root_add_245_5_B_6_,
         add_9_root_add_0_root_add_245_5_B_7_,
         add_9_root_add_0_root_add_245_5_B_8_,
         add_9_root_add_0_root_add_245_5_B_9_,
         add_9_root_add_0_root_add_245_5_B_10_,
         add_9_root_add_0_root_add_245_5_B_11_,
         add_9_root_add_0_root_add_245_5_B_12_,
         add_9_root_add_0_root_add_245_5_B_13_,
         add_9_root_add_0_root_add_245_5_B_14_,
         add_9_root_add_0_root_add_245_5_A_1_,
         add_9_root_add_0_root_add_245_5_A_2_,
         add_9_root_add_0_root_add_245_5_A_3_,
         add_9_root_add_0_root_add_245_5_A_4_,
         add_9_root_add_0_root_add_245_5_A_5_,
         add_9_root_add_0_root_add_245_5_A_6_,
         add_9_root_add_0_root_add_245_5_A_7_,
         add_9_root_add_0_root_add_245_5_A_8_,
         add_9_root_add_0_root_add_245_5_A_9_,
         add_9_root_add_0_root_add_245_5_A_10_,
         add_9_root_add_0_root_add_245_5_A_11_,
         add_9_root_add_0_root_add_245_5_A_12_,
         add_9_root_add_0_root_add_245_5_A_13_,
         add_9_root_add_0_root_add_245_5_A_14_,
         add_9_root_add_0_root_add_245_5_A_15_,
         add_9_root_add_0_root_add_245_5_A_16_,
         add_9_root_add_0_root_add_245_5_A_17_,
         add_9_root_add_0_root_add_245_5_A_18_,
         add_9_root_add_0_root_add_245_5_A_19_,
         add_6_root_add_0_root_add_245_5_carry_5_,
         add_6_root_add_0_root_add_245_5_carry_6_,
         add_6_root_add_0_root_add_245_5_carry_7_,
         add_6_root_add_0_root_add_245_5_carry_8_,
         add_6_root_add_0_root_add_245_5_carry_9_,
         add_6_root_add_0_root_add_245_5_carry_10_,
         add_6_root_add_0_root_add_245_5_carry_11_,
         add_6_root_add_0_root_add_245_5_carry_12_,
         add_6_root_add_0_root_add_245_5_carry_13_,
         add_6_root_add_0_root_add_245_5_carry_14_,
         add_6_root_add_0_root_add_245_5_carry_15_,
         add_6_root_add_0_root_add_245_5_carry_16_,
         add_6_root_add_0_root_add_245_5_carry_17_,
         add_6_root_add_0_root_add_245_5_carry_18_,
         add_6_root_add_0_root_add_245_5_A_3_,
         add_6_root_add_0_root_add_245_5_A_4_,
         add_6_root_add_0_root_add_245_5_A_5_,
         add_6_root_add_0_root_add_245_5_A_6_,
         add_6_root_add_0_root_add_245_5_A_7_,
         add_6_root_add_0_root_add_245_5_A_8_,
         add_6_root_add_0_root_add_245_5_A_9_,
         add_6_root_add_0_root_add_245_5_A_10_,
         add_6_root_add_0_root_add_245_5_A_11_,
         add_6_root_add_0_root_add_245_5_A_12_,
         add_6_root_add_0_root_add_245_5_A_13_,
         add_6_root_add_0_root_add_245_5_A_14_,
         add_6_root_add_0_root_add_245_5_A_15_,
         add_6_root_add_0_root_add_245_5_A_16_,
         add_6_root_add_0_root_add_245_5_A_17_,
         add_7_root_add_0_root_add_245_5_carry_5_,
         add_7_root_add_0_root_add_245_5_carry_6_,
         add_7_root_add_0_root_add_245_5_carry_7_,
         add_7_root_add_0_root_add_245_5_carry_8_,
         add_7_root_add_0_root_add_245_5_carry_9_,
         add_7_root_add_0_root_add_245_5_carry_10_,
         add_7_root_add_0_root_add_245_5_carry_11_,
         add_7_root_add_0_root_add_245_5_carry_12_,
         add_7_root_add_0_root_add_245_5_carry_13_,
         add_7_root_add_0_root_add_245_5_carry_14_,
         add_7_root_add_0_root_add_245_5_carry_15_,
         add_7_root_add_0_root_add_245_5_carry_16_,
         add_7_root_add_0_root_add_245_5_carry_17_,
         add_13_root_add_0_root_add_245_5_carry_5_,
         add_13_root_add_0_root_add_245_5_carry_6_,
         add_13_root_add_0_root_add_245_5_carry_7_,
         add_13_root_add_0_root_add_245_5_carry_8_,
         add_13_root_add_0_root_add_245_5_carry_9_,
         add_13_root_add_0_root_add_245_5_carry_10_,
         add_13_root_add_0_root_add_245_5_carry_11_,
         add_13_root_add_0_root_add_245_5_carry_12_,
         add_13_root_add_0_root_add_245_5_carry_13_,
         add_13_root_add_0_root_add_245_5_carry_14_,
         add_13_root_add_0_root_add_245_5_carry_15_,
         add_13_root_add_0_root_add_245_5_carry_16_,
         add_13_root_add_0_root_add_245_5_carry_17_,
         add_13_root_add_0_root_add_245_5_SUM_3_,
         add_13_root_add_0_root_add_245_5_SUM_4_,
         add_13_root_add_0_root_add_245_5_SUM_5_,
         add_13_root_add_0_root_add_245_5_SUM_6_,
         add_13_root_add_0_root_add_245_5_SUM_7_,
         add_13_root_add_0_root_add_245_5_SUM_8_,
         add_13_root_add_0_root_add_245_5_SUM_9_,
         add_13_root_add_0_root_add_245_5_SUM_10_,
         add_13_root_add_0_root_add_245_5_SUM_11_,
         add_13_root_add_0_root_add_245_5_SUM_12_,
         add_13_root_add_0_root_add_245_5_SUM_13_,
         add_13_root_add_0_root_add_245_5_SUM_14_,
         add_13_root_add_0_root_add_245_5_SUM_15_,
         add_13_root_add_0_root_add_245_5_SUM_16_,
         add_13_root_add_0_root_add_245_5_SUM_17_,
         add_12_root_add_0_root_add_245_5_carry_3_,
         add_12_root_add_0_root_add_245_5_carry_4_,
         add_12_root_add_0_root_add_245_5_carry_5_,
         add_12_root_add_0_root_add_245_5_carry_6_,
         add_12_root_add_0_root_add_245_5_carry_7_,
         add_12_root_add_0_root_add_245_5_carry_8_,
         add_12_root_add_0_root_add_245_5_carry_9_,
         add_12_root_add_0_root_add_245_5_carry_10_,
         add_12_root_add_0_root_add_245_5_carry_11_,
         add_12_root_add_0_root_add_245_5_carry_12_,
         add_12_root_add_0_root_add_245_5_carry_13_,
         add_8_root_add_0_root_add_245_5_carry_5_,
         add_8_root_add_0_root_add_245_5_carry_6_,
         add_8_root_add_0_root_add_245_5_carry_7_,
         add_8_root_add_0_root_add_245_5_carry_8_,
         add_8_root_add_0_root_add_245_5_carry_9_,
         add_8_root_add_0_root_add_245_5_carry_10_,
         add_8_root_add_0_root_add_245_5_carry_11_,
         add_8_root_add_0_root_add_245_5_carry_12_,
         add_8_root_add_0_root_add_245_5_carry_13_,
         add_8_root_add_0_root_add_245_5_carry_14_,
         add_8_root_add_0_root_add_245_5_carry_15_,
         add_8_root_add_0_root_add_245_5_carry_16_, mult_245_5_n23,
         mult_245_5_n22, mult_245_5_n21, mult_245_5_n20, mult_245_5_n19,
         mult_245_5_n18, mult_245_5_n17, mult_245_5_n16, mult_245_5_n15,
         mult_245_5_n14, mult_245_5_n13, mult_245_5_n12, mult_245_5_n11,
         mult_245_5_n10, mult_245_5_n9, mult_245_5_n8, mult_245_5_n7,
         mult_245_5_n6, mult_245_5_n5, mult_245_5_n4, mult_245_5_n3,
         mult_245_5_n2, mult_245_n23, mult_245_n22, mult_245_n21, mult_245_n20,
         mult_245_n19, mult_245_n18, mult_245_n17, mult_245_n16, mult_245_n15,
         mult_245_n14, mult_245_n13, mult_245_n12, mult_245_n11, mult_245_n10,
         mult_245_n9, mult_245_n8, mult_245_n7, mult_245_n6, mult_245_n5,
         mult_245_n4, mult_245_n3, mult_245_n2, mult_244_4_n17, mult_244_4_n16,
         mult_244_4_n15, mult_244_4_n14, mult_244_4_n13, mult_244_4_n12,
         mult_244_4_n11, mult_244_4_n10, mult_244_4_n9, mult_244_4_n8,
         mult_244_4_n7, mult_244_4_n6, mult_244_4_n5, mult_244_4_n4,
         mult_244_4_n3, mult_244_2_n17, mult_244_2_n16, mult_244_2_n15,
         mult_244_2_n14, mult_244_2_n13, mult_244_2_n12, mult_244_2_n11,
         mult_244_2_n10, mult_244_2_n9, mult_244_2_n8, mult_244_2_n7,
         mult_244_2_n6, mult_244_2_n5, mult_244_2_n4, mult_244_2_n3,
         mult_242_4_n17, mult_242_4_n16, mult_242_4_n15, mult_242_4_n14,
         mult_242_4_n13, mult_242_4_n12, mult_242_4_n11, mult_242_4_n10,
         mult_242_4_n9, mult_242_4_n8, mult_242_4_n7, mult_242_4_n6,
         mult_242_4_n5, mult_242_4_n4, mult_242_4_n3, mult_242_2_n17,
         mult_242_2_n16, mult_242_2_n15, mult_242_2_n14, mult_242_2_n13,
         mult_242_2_n12, mult_242_2_n11, mult_242_2_n10, mult_242_2_n9,
         mult_242_2_n8, mult_242_2_n7, mult_242_2_n6, mult_242_2_n5,
         mult_242_2_n4, mult_242_2_n3, mult_241_5_n23, mult_241_5_n22,
         mult_241_5_n21, mult_241_5_n20, mult_241_5_n19, mult_241_5_n18,
         mult_241_5_n17, mult_241_5_n16, mult_241_5_n15, mult_241_5_n14,
         mult_241_5_n13, mult_241_5_n12, mult_241_5_n11, mult_241_5_n10,
         mult_241_5_n9, mult_241_5_n8, mult_241_5_n7, mult_241_5_n6,
         mult_241_5_n5, mult_241_5_n4, mult_241_5_n3, mult_241_5_n2,
         mult_241_n23, mult_241_n22, mult_241_n21, mult_241_n20, mult_241_n19,
         mult_241_n18, mult_241_n17, mult_241_n16, mult_241_n15, mult_241_n14,
         mult_241_n13, mult_241_n12, mult_241_n11, mult_241_n10, mult_241_n9,
         mult_241_n8, mult_241_n7, mult_241_n6, mult_241_n5, mult_241_n4,
         mult_241_n3, mult_241_n2, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n816, n848, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n947, n949, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n9960, n9970, n9980, n9990,
         n10000, n10010, n10020, n10030, n10040, n10050, n10060, n10070,
         n10080, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n12700, n12710, n12720, n12730, n12740, n12750;
  wire   [1:0] state;
  wire   [7:0] row;
  wire   [7:0] col;
  wire   [187:0] array;
  wire   [7:0] i;
  wire   [7:0] j;
  wire   [7:4] add_146_carry;
  wire   [16:2] add_17_root_add_0_root_add_245_5_carry;
  wire   [15:5] add_18_root_add_0_root_add_245_5_carry;
  wire   [15:5] add_19_root_add_0_root_add_245_5_carry;
  wire   [12:3] add_22_root_add_0_root_add_245_5_carry;
  wire   [12:3] add_23_root_add_0_root_add_245_5_carry;
  wire   [15:5] add_20_root_add_0_root_add_245_5_carry;
  wire   [15:5] add_21_root_add_0_root_add_245_5_carry;

  imgproc_DW01_dec_0 sub_257 ( .A({row[6:0], col[6:0]}), .SUM({N2287, N2286, 
        N2285, N2284, N2283, N2282, N2281, N2280, N2279, N2278, N2277, N2276, 
        N2275, N2274}) );
  imgproc_DW01_inc_0 add_236 ( .A(col), .SUM({N1289, N1288, N1287, N1286, 
        N1285, N1284, N1283, N1282}) );
  imgproc_DW01_inc_1 add_225 ( .A(row), .SUM({N1277, N1276, N1275, N1274, 
        N1273, N1272, N1271, N1270}) );
  imgproc_DW01_inc_2 add_151 ( .A({n1290, n1291, n1292, n1293, n1294, n1295, 
        n951, N672, N671, N670, N669, n947, N165, n949}), .SUM({N199, N198, 
        N197, N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186}) );
  imgproc_DW01_inc_3 add_149 ( .A(j), .SUM({N185, N184, N183, N182, N181, N180, 
        N179, N178}) );
  imgproc_DW01_inc_4 r653 ( .A(i), .SUM({N163, N162, N161, N160, N159, N158, 
        N157, N156}) );
  imgproc_DW_mult_uns_23 mult_241_2 ( .a(array[181:174]), .product_15_(N1333), 
        .product_14_(N1332), .product_13_(N1331), .product_12_(N1330), 
        .product_11_(N1329), .product_10_(N1328), .product_9_(N1327), 
        .product_8_(N1326), .product_7_(N1325), .product_6_(N1324), 
        .product_5_(N1323), .product_4_(N1322), .product_3_(N1321) );
  imgproc_DW_mult_uns_22 mult_241_3 ( .a(array[173:166]), .product({N1367, 
        N1366, N1365, N1364, N1363, N1362, N1361, N1360, N1359, N1358, N1357, 
        N1356, N1355, N1354, N1353, N1352, N1351}) );
  imgproc_DW_mult_uns_21 mult_241_4 ( .a(array[165:158]), .product_15_(N1401), 
        .product_14_(N1400), .product_13_(N1399), .product_12_(N1398), 
        .product_11_(N1397), .product_10_(N1396), .product_9_(N1395), 
        .product_8_(N1394), .product_7_(N1393), .product_6_(N1392), 
        .product_5_(N1391), .product_4_(N1390), .product_3_(N1389) );
  imgproc_DW_mult_uns_19 mult_242 ( .a(array[151:144]), .product_15_(N1469), 
        .product_14_(N1468), .product_13_(N1467), .product_12_(N1466), 
        .product_11_(N1465), .product_10_(N1464), .product_9_(N1463), 
        .product_8_(N1462), .product_7_(N1461), .product_6_(N1460), 
        .product_5_(N1459), .product_4_(N1458), .product_3_(N1457) );
  imgproc_DW_mult_uns_17 mult_242_3 ( .a(array[136:129]), .product({N1551, 
        N1550, N1549, N1548, N1547, N1546, N1545, N1544, N1543, N1542, N1541, 
        N1540, N1539, N1538, N1537, N1536, N1535, N1534, N1533, N1532}) );
  imgproc_DW_mult_uns_15 mult_242_5 ( .a(array[121:114]), .product_15_(N1632), 
        .product_14_(N1631), .product_13_(N1630), .product_12_(N1629), 
        .product_11_(N1628), .product_10_(N1627), .product_9_(N1626), 
        .product_8_(N1625), .product_7_(N1624), .product_6_(N1623), 
        .product_5_(N1622), .product_4_(N1621), .product_3_(N1620) );
  imgproc_DW_mult_uns_14 mult_243 ( .a(array[113:106]), .product({N1672, N1671, 
        N1670, N1669, N1668, N1667, N1666, N1665, N1664, N1663, N1662, N1661, 
        N16600, N1659, N1658, N1657, N1656}) );
  imgproc_DW_mult_uns_13 mult_243_2 ( .a(array[105:98]), .product({N1715, 
        N1714, N1713, N1712, N1711, N17100, N1709, N1708, N1707, N1706, N1705, 
        N1704, N1703, N1702, N1701, N17000, N1699, N1698, N1697, N1696}) );
  imgproc_DW_mult_uns_12 mult_243_3 ( .a(array[97:90]), .product_20_(N1759), 
        .product_19_(N1758), .product_18_(N1757), .product_17_(N1756), 
        .product_16_(N1755), .product_15_(N1754), .product_14_(N1753), 
        .product_13_(N1752), .product_12_(N1751), .product_11_(N17500), 
        .product_10_(N1749), .product_9_(N1748), .product_8_(N1747), 
        .product_7_(N1746), .product_6_(N1745), .product_5_(N1744), 
        .product_4_(N1743), .product_3_(N1742) );
  imgproc_DW_mult_uns_11 mult_243_4 ( .a(array[89:82]), .product({N1802, N1801, 
        N18000, N1799, N1798, N1797, N1796, N1795, N1794, N1793, N1792, N1791, 
        N17900, N1789, N1788, N1787, N1786, N1785, N1784, N1783}) );
  imgproc_DW_mult_uns_10 mult_243_5 ( .a(array[81:74]), .product({N1842, N1841, 
        N18400, N1839, N1838, N1837, N1836, N1835, N1834, N1833, N1832, N1831, 
        N18300, N1829, N1828, N1827, N1826}) );
  imgproc_DW_mult_uns_9 mult_244 ( .a(array[73:66]), .product_15_(N1881), 
        .product_14_(N18800), .product_13_(N1879), .product_12_(N1878), 
        .product_11_(N1877), .product_10_(N1876), .product_9_(N1875), 
        .product_8_(N1874), .product_7_(N1873), .product_6_(N1872), 
        .product_5_(N1871), .product_4_(N18700), .product_3_(N1869) );
  imgproc_DW_mult_uns_7 mult_244_3 ( .a(array[58:51]), .product({N1966, N1965, 
        N1964, N1963, N1962, N1961, N19600, N1959, N1958, N1957, N1956, N1955, 
        N1954, N1953, N1952, N1951, N19500, N1949, N1948, N1947}) );
  imgproc_DW_mult_uns_5 mult_244_5 ( .a(array[43:36]), .product_15_(N2047), 
        .product_14_(N2046), .product_13_(N2045), .product_12_(N2044), 
        .product_11_(N2043), .product_10_(N2042), .product_9_(N2041), 
        .product_8_(N2040), .product_7_(N2039), .product_6_(N2038), 
        .product_5_(N2037), .product_4_(N2036), .product_3_(N2035) );
  imgproc_DW_mult_uns_3 mult_245_2 ( .a(array[29:22]), .product_15_(N2122), 
        .product_14_(N2121), .product_13_(N2120), .product_12_(N2119), 
        .product_11_(N2118), .product_10_(N2117), .product_9_(N2116), 
        .product_8_(N2115), .product_7_(N2114), .product_6_(N2113), 
        .product_5_(N2112), .product_4_(N2111), .product_3_(N2110) );
  imgproc_DW_mult_uns_2 mult_245_3 ( .a(array[21:14]), .product({N2162, N2161, 
        N2160, N2159, N2158, N2157, N2156, N2155, N2154, N2153, N2152, N2151, 
        N2150, N2149, N2148, N2147, N2146}) );
  imgproc_DW_mult_uns_1 mult_245_4 ( .a(array[13:6]), .product_15_(N2201), 
        .product_14_(N2200), .product_13_(N2199), .product_12_(N2198), 
        .product_11_(N2197), .product_10_(N2196), .product_9_(N2195), 
        .product_8_(N2194), .product_7_(N2193), .product_6_(N2192), 
        .product_5_(N2191), .product_4_(N2190), .product_3_(N2189) );
  imgproc_DW01_add_19 add_16_root_add_0_root_add_245_5 ( .A_16_(N2162), 
        .A_15_(N2161), .A_14_(N2160), .A_13_(N2159), .A_12_(N2158), .A_11_(
        N2157), .A_10_(N2156), .A_9_(N2155), .A_8_(N2154), .A_7_(N2153), 
        .A_6_(N2152), .A_5_(N2151), .A_4_(N2150), .A_3_(N2149), .A_2_(N2148), 
        .A_1_(N2147), .A_0_(N2146), .B_16_(N1842), .B_15_(N1841), .B_14_(
        N18400), .B_13_(N1839), .B_12_(N1838), .B_11_(N1837), .B_10_(N1836), 
        .B_9_(N1835), .B_8_(N1834), .B_7_(N1833), .B_6_(N1832), .B_5_(N1831), 
        .B_4_(N18300), .B_3_(N1829), .B_2_(N1828), .B_1_(N1827), .B_0_(N1826), 
        .SUM_17_(N1487), .SUM_16_(N1486), .SUM_15_(N1485), .SUM_14_(N1484), 
        .SUM_13_(N1483), .SUM_12_(N1482), .SUM_11_(N1481), .SUM_10_(N1480), 
        .SUM_9_(N1479), .SUM_8_(N1478), .SUM_7_(N1477), .SUM_6_(N1476), 
        .SUM_5_(N1475), .SUM_4_(N1474), .SUM_3_(N1473), .SUM_2_(N1472), 
        .SUM_1_(N1471), .SUM_0_(N1470) );
  imgproc_DW01_add_16 add_15_root_add_0_root_add_245_5 ( .A_18_(N1593), 
        .A_17_(N1592), .A_16_(N1591), .A_15_(N1590), .A_14_(N1589), .A_13_(
        N1588), .A_12_(N1587), .A_11_(N1586), .A_10_(N1585), .A_9_(N1584), 
        .A_8_(N1583), .A_7_(N1582), .A_6_(N1581), .A_5_(N1580), .A_4_(N1579), 
        .A_3_(N1578), .A_2_(N1577), .A_1_(N1576), .A_0_(N1575), .B_18_(N2008), 
        .B_17_(N2007), .B_16_(N2006), .B_15_(N2005), .B_14_(N2004), .B_13_(
        N2003), .B_12_(N2002), .B_11_(N2001), .B_10_(N2000), .B_9_(N1999), 
        .B_8_(N1998), .B_7_(N1997), .B_6_(N1996), .B_5_(N1995), .B_4_(N1994), 
        .B_3_(N1993), .B_2_(N1992), .B_1_(N1991), .B_0_(N19900), .SUM_19_(
        add_9_root_add_0_root_add_245_5_A_19_), .SUM_18_(
        add_9_root_add_0_root_add_245_5_A_18_), .SUM_17_(
        add_9_root_add_0_root_add_245_5_A_17_), .SUM_16_(
        add_9_root_add_0_root_add_245_5_A_16_), .SUM_15_(
        add_9_root_add_0_root_add_245_5_A_15_), .SUM_14_(
        add_9_root_add_0_root_add_245_5_A_14_), .SUM_13_(
        add_9_root_add_0_root_add_245_5_A_13_), .SUM_12_(
        add_9_root_add_0_root_add_245_5_A_12_), .SUM_11_(
        add_9_root_add_0_root_add_245_5_A_11_), .SUM_10_(
        add_9_root_add_0_root_add_245_5_A_10_), .SUM_9_(
        add_9_root_add_0_root_add_245_5_A_9_), .SUM_8_(
        add_9_root_add_0_root_add_245_5_A_8_), .SUM_7_(
        add_9_root_add_0_root_add_245_5_A_7_), .SUM_6_(
        add_9_root_add_0_root_add_245_5_A_6_), .SUM_5_(
        add_9_root_add_0_root_add_245_5_A_5_), .SUM_4_(
        add_9_root_add_0_root_add_245_5_A_4_), .SUM_3_(
        add_9_root_add_0_root_add_245_5_A_3_), .SUM_2_(
        add_9_root_add_0_root_add_245_5_A_2_), .SUM_1_(
        add_9_root_add_0_root_add_245_5_A_1_), .SUM_0_(N2202) );
  imgproc_DW01_add_15 add_11_root_add_0_root_add_245_5 ( .A_19_(N1802), 
        .A_18_(N1801), .A_17_(N18000), .A_16_(N1799), .A_15_(N1798), .A_14_(
        N1797), .A_13_(N1796), .A_12_(N1795), .A_11_(N1794), .A_10_(N1793), 
        .A_9_(N1792), .A_8_(N1791), .A_7_(N17900), .A_6_(N1789), .A_5_(N1788), 
        .A_4_(N1787), .A_3_(N1786), .A_2_(N1785), .A_1_(N1784), .A_0_(N1783), 
        .B_19_(N1715), .B_18_(N1714), .B_17_(N1713), .B_16_(N1712), .B_15_(
        N1711), .B_14_(N17100), .B_13_(N1709), .B_12_(N1708), .B_11_(N1707), 
        .B_10_(N1706), .B_9_(N1705), .B_8_(N1704), .B_7_(N1703), .B_6_(N1702), 
        .B_5_(N1701), .B_4_(N17000), .B_3_(N1699), .B_2_(N1698), .B_1_(N1697), 
        .B_0_(N1696), .SUM_20_(N1863), .SUM_19_(N1862), .SUM_18_(N1861), 
        .SUM_17_(N18600), .SUM_16_(N1859), .SUM_15_(N1858), .SUM_14_(N1857), 
        .SUM_13_(N1856), .SUM_12_(N1855), .SUM_11_(N1854), .SUM_10_(N1853), 
        .SUM_9_(N1852), .SUM_8_(N1851), .SUM_7_(N18500), .SUM_6_(N1849), 
        .SUM_5_(N1848), .SUM_4_(N1847), .SUM_3_(N1846), .SUM_2_(N1845), 
        .SUM_1_(N1844), .SUM_0_(N1843) );
  imgproc_DW01_add_14 add_10_root_add_0_root_add_245_5 ( .A_19_(N1551), 
        .A_18_(N1550), .A_17_(N1549), .A_16_(N1548), .A_15_(N1547), .A_14_(
        N1546), .A_13_(N1545), .A_12_(N1544), .A_11_(N1543), .A_10_(N1542), 
        .A_9_(N1541), .A_8_(N1540), .A_7_(N1539), .A_6_(N1538), .A_5_(N1537), 
        .A_4_(N1536), .A_3_(N1535), .A_2_(N1534), .A_1_(N1533), .A_0_(N1532), 
        .B_19_(N1966), .B_18_(N1965), .B_17_(N1964), .B_16_(N1963), .B_15_(
        N1962), .B_14_(N1961), .B_13_(N19600), .B_12_(N1959), .B_11_(N1958), 
        .B_10_(N1957), .B_9_(N1956), .B_8_(N1955), .B_7_(N1954), .B_6_(N1953), 
        .B_5_(N1952), .B_4_(N1951), .B_3_(N19500), .B_2_(N1949), .B_1_(N1948), 
        .B_0_(N1947), .SUM_20_(N2104), .SUM_19_(N2103), .SUM_18_(N2102), 
        .SUM_17_(N2101), .SUM_16_(N2100), .SUM_15_(N2099), .SUM_14_(N2098), 
        .SUM_13_(N2097), .SUM_12_(N2096), .SUM_11_(N2095), .SUM_10_(N2094), 
        .SUM_9_(N2093), .SUM_8_(N2092), .SUM_7_(N2091), .SUM_6_(N2090), 
        .SUM_5_(N2089), .SUM_4_(N2088), .SUM_3_(N2087), .SUM_2_(N2086), 
        .SUM_1_(N2085), .SUM_0_(N2084) );
  imgproc_DW01_add_13 add_3_root_add_0_root_add_245_5 ( .A_20_(N1863), .A_19_(
        N1862), .A_18_(N1861), .A_17_(N18600), .A_16_(N1859), .A_15_(N1858), 
        .A_14_(N1857), .A_13_(N1856), .A_12_(N1855), .A_11_(N1854), .A_10_(
        N1853), .A_9_(N1852), .A_8_(N1851), .A_7_(N18500), .A_6_(N1849), 
        .A_5_(N1848), .A_4_(N1847), .A_3_(N1846), .A_2_(N1845), .A_1_(N1844), 
        .A_0_(N1843), .B_20_(N2104), .B_19_(N2103), .B_18_(N2102), .B_17_(
        N2101), .B_16_(N2100), .B_15_(N2099), .B_14_(N2098), .B_13_(N2097), 
        .B_12_(N2096), .B_11_(N2095), .B_10_(N2094), .B_9_(N2093), .B_8_(N2092), .B_7_(N2091), .B_6_(N2090), .B_5_(N2089), .B_4_(N2088), .B_3_(N2087), .B_2_(
        N2086), .B_1_(N2085), .B_0_(N2084), .SUM_21_(N1694), .SUM_20_(N1693), 
        .SUM_19_(N1692), .SUM_18_(N1691), .SUM_17_(N16900), .SUM_16_(N1689), 
        .SUM_15_(N1688), .SUM_14_(N1687), .SUM_13_(N1686), .SUM_12_(N1685), 
        .SUM_11_(N1684), .SUM_10_(N1683), .SUM_9_(N1682), .SUM_8_(N1681), 
        .SUM_7_(N16800), .SUM_6_(N1679), .SUM_5_(N1678), .SUM_4_(N1677), 
        .SUM_3_(N1676), .SUM_2_(N1675), .SUM_1_(N1674), .SUM_0_(N1673) );
  imgproc_DW01_add_9 add_5_root_add_0_root_add_245_5 ( .A_18_(n806), .A_17_(
        N18200), .A_16_(N1819), .A_15_(N1818), .A_14_(N1817), .A_13_(N1816), 
        .A_12_(N1815), .A_11_(N1814), .A_10_(N1813), .A_9_(N1812), .A_8_(N1811), .A_7_(N18100), .A_6_(N1809), .A_5_(N1808), .A_4_(N1807), .A_3_(N1806), 
        .A_2_(N1805), .A_1_(N1804), .A_0_(N1803), .B_18_(n794), .B_17_(
        add_13_root_add_0_root_add_245_5_SUM_17_), .B_16_(
        add_13_root_add_0_root_add_245_5_SUM_16_), .B_15_(
        add_13_root_add_0_root_add_245_5_SUM_15_), .B_14_(
        add_13_root_add_0_root_add_245_5_SUM_14_), .B_13_(
        add_13_root_add_0_root_add_245_5_SUM_13_), .B_12_(
        add_13_root_add_0_root_add_245_5_SUM_12_), .B_11_(
        add_13_root_add_0_root_add_245_5_SUM_11_), .B_10_(
        add_13_root_add_0_root_add_245_5_SUM_10_), .B_9_(
        add_13_root_add_0_root_add_245_5_SUM_9_), .B_8_(
        add_13_root_add_0_root_add_245_5_SUM_8_), .B_7_(
        add_13_root_add_0_root_add_245_5_SUM_7_), .B_6_(
        add_13_root_add_0_root_add_245_5_SUM_6_), .B_5_(
        add_13_root_add_0_root_add_245_5_SUM_5_), .B_4_(
        add_13_root_add_0_root_add_245_5_SUM_4_), .B_3_(
        add_13_root_add_0_root_add_245_5_SUM_3_), .B_2_(N1472), .B_1_(N1471), 
        .B_0_(N1470), .SUM_19_(N2067), .SUM_18_(N2066), .SUM_17_(N2065), 
        .SUM_16_(N2064), .SUM_15_(N2063), .SUM_14_(N2062), .SUM_13_(N2061), 
        .SUM_12_(N2060), .SUM_11_(N2059), .SUM_10_(N2058), .SUM_9_(N2057), 
        .SUM_8_(N2056), .SUM_7_(N2055), .SUM_6_(N2054), .SUM_5_(N2053), 
        .SUM_4_(N2052), .SUM_3_(N2051), .SUM_2_(N2050), .SUM_1_(N2049), 
        .SUM_0_(N2048) );
  imgproc_DW01_add_8 add_14_root_add_0_root_add_245_5 ( .A_18_(N1509), .A_17_(
        N1508), .A_16_(N1507), .A_15_(N1506), .A_14_(N1505), .A_13_(N1504), 
        .A_12_(N1503), .A_11_(N1502), .A_10_(N1501), .A_9_(N1500), .A_8_(N1499), .A_7_(N1498), .A_6_(N1497), .A_5_(N1496), .A_4_(N1495), .A_3_(N1494), .A_2_(
        N1493), .A_1_(N1492), .A_0_(N1491), .B_18_(N1923), .B_17_(N1922), 
        .B_16_(N1921), .B_15_(N19200), .B_14_(N1919), .B_13_(N1918), .B_12_(
        N1917), .B_11_(N1916), .B_10_(N1915), .B_9_(N1914), .B_8_(N1913), 
        .B_7_(N1912), .B_6_(N1911), .B_5_(N19100), .B_4_(N1909), .B_3_(N1908), 
        .B_2_(N1907), .B_1_(N1906), .B_0_(N1905), .SUM_19_(N1901), .SUM_18_(
        N19000), .SUM_17_(N1899), .SUM_16_(N1898), .SUM_15_(N1897), .SUM_14_(
        N1896), .SUM_13_(N1895), .SUM_12_(N1894), .SUM_11_(N1893), .SUM_10_(
        N1892), .SUM_9_(N1891), .SUM_8_(N18900), .SUM_7_(N1889), .SUM_6_(N1888), .SUM_5_(N1887), .SUM_4_(N1886), .SUM_3_(N1885), .SUM_2_(N1884), .SUM_1_(
        N1883), .SUM_0_(N1882) );
  imgproc_DW01_add_7 add_4_root_add_0_root_add_245_5 ( .A_19_(N2067), .A_18_(
        N2066), .A_17_(N2065), .A_16_(N2064), .A_15_(N2063), .A_14_(N2062), 
        .A_13_(N2061), .A_12_(N2060), .A_11_(N2059), .A_10_(N2058), .A_9_(
        N2057), .A_8_(N2056), .A_7_(N2055), .A_6_(N2054), .A_5_(N2053), .A_4_(
        N2052), .A_3_(N2051), .A_2_(N2050), .A_1_(N2049), .A_0_(N2048), 
        .B_19_(N1901), .B_18_(N19000), .B_17_(N1899), .B_16_(N1898), .B_15_(
        N1897), .B_14_(N1896), .B_13_(N1895), .B_12_(N1894), .B_11_(N1893), 
        .B_10_(N1892), .B_9_(N1891), .B_8_(N18900), .B_7_(N1889), .B_6_(N1888), 
        .B_5_(N1887), .B_4_(N1886), .B_3_(N1885), .B_2_(N1884), .B_1_(N1883), 
        .B_0_(N1882), .SUM_20_(N1736), .SUM_19_(N1735), .SUM_18_(N1734), 
        .SUM_17_(N1733), .SUM_16_(N1732), .SUM_15_(N1731), .SUM_14_(N17300), 
        .SUM_13_(N1729), .SUM_12_(N1728), .SUM_11_(N1727), .SUM_10_(N1726), 
        .SUM_9_(N1725), .SUM_8_(N1724), .SUM_7_(N1723), .SUM_6_(N1722), 
        .SUM_5_(N1721), .SUM_4_(N17200), .SUM_3_(N1719), .SUM_2_(N1718), 
        .SUM_1_(N1717), .SUM_0_(N1716) );
  imgproc_DW01_add_4 add_2_root_add_0_root_add_245_5 ( .A_20_(N1736), .A_19_(
        N1735), .A_18_(N1734), .A_17_(N1733), .A_16_(N1732), .A_15_(N1731), 
        .A_14_(N17300), .A_13_(N1729), .A_12_(N1728), .A_11_(N1727), .A_10_(
        N1726), .A_9_(N1725), .A_8_(N1724), .A_7_(N1723), .A_6_(N1722), .A_5_(
        N1721), .A_4_(N17200), .A_3_(N1719), .A_2_(N1718), .A_1_(N1717), 
        .A_0_(N1716), .B_20_(n811), .B_19_(N2221), .B_18_(N2220), .B_17_(N2219), .B_16_(N2218), .B_15_(N2217), .B_14_(N2216), .B_13_(N2215), .B_12_(N2214), 
        .B_11_(N2213), .B_10_(N2212), .B_9_(N2211), .B_8_(N2210), .B_7_(N2209), 
        .B_6_(N2208), .B_5_(N2207), .B_4_(N2206), .B_3_(N2205), .B_2_(N2204), 
        .B_1_(N2203), .B_0_(N2202), .SUM_21_(N2030), .SUM_20_(N2029), 
        .SUM_19_(N2028), .SUM_18_(N2027), .SUM_17_(N2026), .SUM_16_(N2025), 
        .SUM_15_(N2024), .SUM_14_(N2023), .SUM_13_(N2022), .SUM_12_(N2021), 
        .SUM_11_(N2020), .SUM_10_(N2019), .SUM_9_(N2018), .SUM_8_(N2017), 
        .SUM_7_(N2016), .SUM_6_(N2015), .SUM_5_(N2014), .SUM_4_(N2013), 
        .SUM_3_(N2012), .SUM_2_(N2011), .SUM_1_(N2010), .SUM_0_(N2009) );
  imgproc_DW01_add_3 add_1_root_add_0_root_add_245_5 ( .SUM({N2185, N2184, 
        N2183, N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, 
        N2173, N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, 
        N2163}), .A_21_(n812), .A_20_(N17800), .A_19_(N1779), .A_18_(N1778), 
        .A_17_(N1777), .A_16_(N1776), .A_15_(N1775), .A_14_(N1774), .A_13_(
        N1773), .A_12_(N1772), .A_11_(N1771), .A_10_(N17700), .A_9_(N1769), 
        .A_8_(N1768), .A_7_(N1767), .A_6_(N1766), .A_5_(N1765), .A_4_(N1764), 
        .A_3_(N1763), .B_21_(N1694), .B_20_(N1693), .B_19_(N1692), .B_18_(
        N1691), .B_17_(N16900), .B_16_(N1689), .B_15_(N1688), .B_14_(N1687), 
        .B_13_(N1686), .B_12_(N1685), .B_11_(N1684), .B_10_(N1683), .B_9_(
        N1682), .B_8_(N1681), .B_7_(N16800), .B_6_(N1679), .B_5_(N1678), 
        .B_4_(N1677), .B_3_(N1676), .B_2_(N1675), .B_1_(N1674), .B_0_(N1673)
         );
  imgproc_DW01_add_2 add_0_root_add_0_root_add_245_5 ( .B({N2185, N2184, N2183, 
        N2182, N2181, N2180, N2179, N2178, N2177, N2176, N2175, N2174, N2173, 
        N2172, N2171, N2170, N2169, N2168, N2167, N2166, N2165, N2164, N2163}), 
        .A_21_(N2030), .A_20_(N2029), .A_19_(N2028), .A_18_(N2027), .A_17_(
        N2026), .A_16_(N2025), .A_15_(N2024), .A_14_(N2023), .A_13_(N2022), 
        .A_12_(N2021), .A_11_(N2020), .A_10_(N2019), .A_9_(N2018), .A_8_(N2017), .A_7_(N2016), .A_6_(N2015), .A_5_(N2014), .A_4_(N2013), .A_3_(N2012), .A_2_(
        N2011), .A_1_(N2010), .A_0_(N2009), .SUM_22_(N2246), .SUM_21_(N2245), 
        .SUM_20_(N2244), .SUM_19_(N2243), .SUM_18_(N2242), .SUM_17_(N2241), 
        .SUM_16_(N2240), .SUM_15_(N2239), .SUM_14_(N2238) );
  imgproc_DW01_inc_5 add_250 ( .A({N2246, n792, N2244, N2243, N2242, N2241, 
        N2240, N2239}), .SUM({N2257, N2256, N2255, N2254, N2253, N2252, N2251, 
        N2250}) );
  ADDHXL mult_245_5_U17 ( .A(array[1]), .B(N2227), .CO(mult_245_5_n22), .S(
        mult_245_5_n23) );
  ADDFXL mult_245_5_U16 ( .A(N2227), .B(array[2]), .CI(array[0]), .CO(
        mult_245_5_n20), .S(mult_245_5_n21) );
  ADDFXL mult_245_5_U15 ( .A(array[0]), .B(array[3]), .CI(array[1]), .CO(
        mult_245_5_n18), .S(mult_245_5_n19) );
  ADDFXL mult_245_5_U14 ( .A(array[1]), .B(array[4]), .CI(array[2]), .CO(
        mult_245_5_n16), .S(mult_245_5_n17) );
  ADDFXL mult_245_5_U13 ( .A(array[2]), .B(array[5]), .CI(array[3]), .CO(
        mult_245_5_n14), .S(mult_245_5_n15) );
  ADDHXL mult_245_5_U12 ( .A(array[4]), .B(array[3]), .CO(mult_245_5_n12), .S(
        mult_245_5_n13) );
  ADDHXL mult_245_5_U11 ( .A(array[5]), .B(array[4]), .CO(mult_245_5_n10), .S(
        mult_245_5_n11) );
  ADDHXL mult_245_5_U10 ( .A(N2226), .B(array[0]), .CO(mult_245_5_n9), .S(
        N2228) );
  ADDFXL mult_245_5_U9 ( .A(mult_245_5_n9), .B(N2226), .CI(mult_245_5_n23), 
        .CO(mult_245_5_n8), .S(N2229) );
  ADDFXL mult_245_5_U8 ( .A(mult_245_5_n21), .B(mult_245_5_n22), .CI(
        mult_245_5_n8), .CO(mult_245_5_n7), .S(N2230) );
  ADDFXL mult_245_5_U7 ( .A(mult_245_5_n19), .B(mult_245_5_n20), .CI(
        mult_245_5_n7), .CO(mult_245_5_n6), .S(N2231) );
  ADDFXL mult_245_5_U6 ( .A(mult_245_5_n17), .B(mult_245_5_n18), .CI(
        mult_245_5_n6), .CO(mult_245_5_n5), .S(N2232) );
  ADDFXL mult_245_5_U5 ( .A(mult_245_5_n15), .B(mult_245_5_n16), .CI(
        mult_245_5_n5), .CO(mult_245_5_n4), .S(N2233) );
  ADDFXL mult_245_5_U4 ( .A(mult_245_5_n14), .B(mult_245_5_n13), .CI(
        mult_245_5_n4), .CO(mult_245_5_n3), .S(N2234) );
  ADDFXL mult_245_5_U3 ( .A(mult_245_5_n11), .B(mult_245_5_n12), .CI(
        mult_245_5_n3), .CO(mult_245_5_n2), .S(N2235) );
  ADDFXL mult_245_5_U2 ( .A(mult_245_5_n10), .B(array[5]), .CI(mult_245_5_n2), 
        .CO(N2237), .S(N2236) );
  ADDHXL mult_245_U17 ( .A(array[31]), .B(N2073), .CO(mult_245_n22), .S(
        mult_245_n23) );
  ADDFXL mult_245_U16 ( .A(N2073), .B(array[32]), .CI(array[30]), .CO(
        mult_245_n20), .S(mult_245_n21) );
  ADDFXL mult_245_U15 ( .A(array[30]), .B(array[33]), .CI(array[31]), .CO(
        mult_245_n18), .S(mult_245_n19) );
  ADDFXL mult_245_U14 ( .A(array[31]), .B(array[34]), .CI(array[32]), .CO(
        mult_245_n16), .S(mult_245_n17) );
  ADDFXL mult_245_U13 ( .A(array[32]), .B(array[35]), .CI(array[33]), .CO(
        mult_245_n14), .S(mult_245_n15) );
  ADDHXL mult_245_U12 ( .A(array[34]), .B(array[33]), .CO(mult_245_n12), .S(
        mult_245_n13) );
  ADDHXL mult_245_U11 ( .A(array[35]), .B(array[34]), .CO(mult_245_n10), .S(
        mult_245_n11) );
  ADDHXL mult_245_U10 ( .A(N2072), .B(array[30]), .CO(mult_245_n9), .S(N2074)
         );
  ADDFXL mult_245_U9 ( .A(mult_245_n9), .B(N2072), .CI(mult_245_n23), .CO(
        mult_245_n8), .S(N2075) );
  ADDFXL mult_245_U8 ( .A(mult_245_n21), .B(mult_245_n22), .CI(mult_245_n8), 
        .CO(mult_245_n7), .S(N2076) );
  ADDFXL mult_245_U7 ( .A(mult_245_n19), .B(mult_245_n20), .CI(mult_245_n7), 
        .CO(mult_245_n6), .S(N2077) );
  ADDFXL mult_245_U6 ( .A(mult_245_n17), .B(mult_245_n18), .CI(mult_245_n6), 
        .CO(mult_245_n5), .S(N2078) );
  ADDFXL mult_245_U5 ( .A(mult_245_n15), .B(mult_245_n16), .CI(mult_245_n5), 
        .CO(mult_245_n4), .S(N2079) );
  ADDFXL mult_245_U4 ( .A(mult_245_n14), .B(mult_245_n13), .CI(mult_245_n4), 
        .CO(mult_245_n3), .S(N2080) );
  ADDFXL mult_245_U3 ( .A(mult_245_n11), .B(mult_245_n12), .CI(mult_245_n3), 
        .CO(mult_245_n2), .S(N2081) );
  ADDFXL mult_245_U2 ( .A(mult_245_n10), .B(array[35]), .CI(mult_245_n2), .CO(
        N2083), .S(N2082) );
  ADDHXL mult_244_4_U20 ( .A(n10050), .B(n10040), .CO(mult_244_4_n17), .S(
        N1991) );
  ADDHXL mult_244_4_U19 ( .A(n10060), .B(mult_244_4_n17), .CO(mult_244_4_n16), 
        .S(N1992) );
  ADDFXL mult_244_4_U18 ( .A(N19900), .B(n10070), .CI(mult_244_4_n16), .CO(
        mult_244_4_n15), .S(N1993) );
  ADDFXL mult_244_4_U17 ( .A(array[44]), .B(n10080), .CI(mult_244_4_n15), .CO(
        mult_244_4_n14), .S(N1994) );
  ADDFXL mult_244_4_U16 ( .A(array[45]), .B(n1009), .CI(mult_244_4_n14), .CO(
        mult_244_4_n13), .S(N1995) );
  ADDFXL mult_244_4_U15 ( .A(array[46]), .B(n1010), .CI(mult_244_4_n13), .CO(
        mult_244_4_n12), .S(N1996) );
  ADDFXL mult_244_4_U14 ( .A(array[47]), .B(n1011), .CI(mult_244_4_n12), .CO(
        mult_244_4_n11), .S(N1997) );
  ADDFXL mult_244_4_U13 ( .A(array[48]), .B(n10040), .CI(mult_244_4_n11), .CO(
        mult_244_4_n10), .S(N1998) );
  ADDFXL mult_244_4_U12 ( .A(array[49]), .B(n10050), .CI(mult_244_4_n10), .CO(
        mult_244_4_n9), .S(N1999) );
  ADDFXL mult_244_4_U11 ( .A(array[50]), .B(n10060), .CI(mult_244_4_n9), .CO(
        mult_244_4_n8), .S(N2000) );
  ADDFXL mult_244_4_U10 ( .A(N19900), .B(n10070), .CI(mult_244_4_n8), .CO(
        mult_244_4_n7), .S(N2001) );
  ADDFXL mult_244_4_U9 ( .A(array[44]), .B(n10080), .CI(mult_244_4_n7), .CO(
        mult_244_4_n6), .S(N2002) );
  ADDFXL mult_244_4_U8 ( .A(array[45]), .B(n1009), .CI(mult_244_4_n6), .CO(
        mult_244_4_n5), .S(N2003) );
  ADDFXL mult_244_4_U7 ( .A(array[46]), .B(n1010), .CI(mult_244_4_n5), .CO(
        mult_244_4_n4), .S(N2004) );
  ADDFXL mult_244_4_U6 ( .A(array[47]), .B(n1011), .CI(mult_244_4_n4), .CO(
        mult_244_4_n3), .S(N2005) );
  ADDHXL mult_244_2_U20 ( .A(n995), .B(n994), .CO(mult_244_2_n17), .S(N1906)
         );
  ADDHXL mult_244_2_U19 ( .A(n9960), .B(mult_244_2_n17), .CO(mult_244_2_n16), 
        .S(N1907) );
  ADDFXL mult_244_2_U18 ( .A(N1905), .B(n9970), .CI(mult_244_2_n16), .CO(
        mult_244_2_n15), .S(N1908) );
  ADDFXL mult_244_2_U17 ( .A(array[59]), .B(n9980), .CI(mult_244_2_n15), .CO(
        mult_244_2_n14), .S(N1909) );
  ADDFXL mult_244_2_U16 ( .A(array[60]), .B(n9990), .CI(mult_244_2_n14), .CO(
        mult_244_2_n13), .S(N19100) );
  ADDFXL mult_244_2_U15 ( .A(array[61]), .B(n10000), .CI(mult_244_2_n13), .CO(
        mult_244_2_n12), .S(N1911) );
  ADDFXL mult_244_2_U14 ( .A(array[62]), .B(n10010), .CI(mult_244_2_n12), .CO(
        mult_244_2_n11), .S(N1912) );
  ADDFXL mult_244_2_U13 ( .A(array[63]), .B(n994), .CI(mult_244_2_n11), .CO(
        mult_244_2_n10), .S(N1913) );
  ADDFXL mult_244_2_U12 ( .A(array[64]), .B(n995), .CI(mult_244_2_n10), .CO(
        mult_244_2_n9), .S(N1914) );
  ADDFXL mult_244_2_U11 ( .A(array[65]), .B(n9960), .CI(mult_244_2_n9), .CO(
        mult_244_2_n8), .S(N1915) );
  ADDFXL mult_244_2_U10 ( .A(N1905), .B(n9970), .CI(mult_244_2_n8), .CO(
        mult_244_2_n7), .S(N1916) );
  ADDFXL mult_244_2_U9 ( .A(array[59]), .B(n9980), .CI(mult_244_2_n7), .CO(
        mult_244_2_n6), .S(N1917) );
  ADDFXL mult_244_2_U8 ( .A(array[60]), .B(n9990), .CI(mult_244_2_n6), .CO(
        mult_244_2_n5), .S(N1918) );
  ADDFXL mult_244_2_U7 ( .A(array[61]), .B(n10000), .CI(mult_244_2_n5), .CO(
        mult_244_2_n4), .S(N1919) );
  ADDFXL mult_244_2_U6 ( .A(array[62]), .B(n10010), .CI(mult_244_2_n4), .CO(
        mult_244_2_n3), .S(N19200) );
  ADDHXL mult_242_4_U20 ( .A(n985), .B(n984), .CO(mult_242_4_n17), .S(N1576)
         );
  ADDHXL mult_242_4_U19 ( .A(n986), .B(mult_242_4_n17), .CO(mult_242_4_n16), 
        .S(N1577) );
  ADDFXL mult_242_4_U18 ( .A(N1575), .B(n987), .CI(mult_242_4_n16), .CO(
        mult_242_4_n15), .S(N1578) );
  ADDFXL mult_242_4_U17 ( .A(array[122]), .B(n988), .CI(mult_242_4_n15), .CO(
        mult_242_4_n14), .S(N1579) );
  ADDFXL mult_242_4_U16 ( .A(array[123]), .B(n989), .CI(mult_242_4_n14), .CO(
        mult_242_4_n13), .S(N1580) );
  ADDFXL mult_242_4_U15 ( .A(array[124]), .B(n990), .CI(mult_242_4_n13), .CO(
        mult_242_4_n12), .S(N1581) );
  ADDFXL mult_242_4_U14 ( .A(array[125]), .B(n991), .CI(mult_242_4_n12), .CO(
        mult_242_4_n11), .S(N1582) );
  ADDFXL mult_242_4_U13 ( .A(array[126]), .B(n984), .CI(mult_242_4_n11), .CO(
        mult_242_4_n10), .S(N1583) );
  ADDFXL mult_242_4_U12 ( .A(array[127]), .B(n985), .CI(mult_242_4_n10), .CO(
        mult_242_4_n9), .S(N1584) );
  ADDFXL mult_242_4_U11 ( .A(array[128]), .B(n986), .CI(mult_242_4_n9), .CO(
        mult_242_4_n8), .S(N1585) );
  ADDFXL mult_242_4_U10 ( .A(N1575), .B(n987), .CI(mult_242_4_n8), .CO(
        mult_242_4_n7), .S(N1586) );
  ADDFXL mult_242_4_U9 ( .A(array[122]), .B(n988), .CI(mult_242_4_n7), .CO(
        mult_242_4_n6), .S(N1587) );
  ADDFXL mult_242_4_U8 ( .A(array[123]), .B(n989), .CI(mult_242_4_n6), .CO(
        mult_242_4_n5), .S(N1588) );
  ADDFXL mult_242_4_U7 ( .A(array[124]), .B(n990), .CI(mult_242_4_n5), .CO(
        mult_242_4_n4), .S(N1589) );
  ADDFXL mult_242_4_U6 ( .A(array[125]), .B(n991), .CI(mult_242_4_n4), .CO(
        mult_242_4_n3), .S(N1590) );
  ADDHXL mult_242_2_U20 ( .A(n975), .B(n974), .CO(mult_242_2_n17), .S(N1492)
         );
  ADDHXL mult_242_2_U19 ( .A(n976), .B(mult_242_2_n17), .CO(mult_242_2_n16), 
        .S(N1493) );
  ADDFXL mult_242_2_U18 ( .A(N1491), .B(n977), .CI(mult_242_2_n16), .CO(
        mult_242_2_n15), .S(N1494) );
  ADDFXL mult_242_2_U17 ( .A(array[137]), .B(n978), .CI(mult_242_2_n15), .CO(
        mult_242_2_n14), .S(N1495) );
  ADDFXL mult_242_2_U16 ( .A(array[138]), .B(n979), .CI(mult_242_2_n14), .CO(
        mult_242_2_n13), .S(N1496) );
  ADDFXL mult_242_2_U15 ( .A(array[139]), .B(n980), .CI(mult_242_2_n13), .CO(
        mult_242_2_n12), .S(N1497) );
  ADDFXL mult_242_2_U14 ( .A(array[140]), .B(n981), .CI(mult_242_2_n12), .CO(
        mult_242_2_n11), .S(N1498) );
  ADDFXL mult_242_2_U13 ( .A(array[141]), .B(n974), .CI(mult_242_2_n11), .CO(
        mult_242_2_n10), .S(N1499) );
  ADDFXL mult_242_2_U12 ( .A(array[142]), .B(n975), .CI(mult_242_2_n10), .CO(
        mult_242_2_n9), .S(N1500) );
  ADDFXL mult_242_2_U11 ( .A(array[143]), .B(n976), .CI(mult_242_2_n9), .CO(
        mult_242_2_n8), .S(N1501) );
  ADDFXL mult_242_2_U10 ( .A(N1491), .B(n977), .CI(mult_242_2_n8), .CO(
        mult_242_2_n7), .S(N1502) );
  ADDFXL mult_242_2_U9 ( .A(array[137]), .B(n978), .CI(mult_242_2_n7), .CO(
        mult_242_2_n6), .S(N1503) );
  ADDFXL mult_242_2_U8 ( .A(array[138]), .B(n979), .CI(mult_242_2_n6), .CO(
        mult_242_2_n5), .S(N1504) );
  ADDFXL mult_242_2_U7 ( .A(array[139]), .B(n980), .CI(mult_242_2_n5), .CO(
        mult_242_2_n4), .S(N1505) );
  ADDFXL mult_242_2_U6 ( .A(array[140]), .B(n981), .CI(mult_242_2_n4), .CO(
        mult_242_2_n3), .S(N1506) );
  ADDHXL mult_241_5_U17 ( .A(array[153]), .B(N1423), .CO(mult_241_5_n22), .S(
        mult_241_5_n23) );
  ADDFXL mult_241_5_U16 ( .A(N1423), .B(array[154]), .CI(array[152]), .CO(
        mult_241_5_n20), .S(mult_241_5_n21) );
  ADDFXL mult_241_5_U15 ( .A(array[152]), .B(array[155]), .CI(array[153]), 
        .CO(mult_241_5_n18), .S(mult_241_5_n19) );
  ADDFXL mult_241_5_U14 ( .A(array[153]), .B(array[156]), .CI(array[154]), 
        .CO(mult_241_5_n16), .S(mult_241_5_n17) );
  ADDFXL mult_241_5_U13 ( .A(array[154]), .B(array[157]), .CI(array[155]), 
        .CO(mult_241_5_n14), .S(mult_241_5_n15) );
  ADDHXL mult_241_5_U12 ( .A(array[156]), .B(array[155]), .CO(mult_241_5_n12), 
        .S(mult_241_5_n13) );
  ADDHXL mult_241_5_U11 ( .A(array[157]), .B(array[156]), .CO(mult_241_5_n10), 
        .S(mult_241_5_n11) );
  ADDHXL mult_241_5_U10 ( .A(N1422), .B(array[152]), .CO(mult_241_5_n9), .S(
        N1424) );
  ADDFXL mult_241_5_U9 ( .A(mult_241_5_n9), .B(N1422), .CI(mult_241_5_n23), 
        .CO(mult_241_5_n8), .S(N1425) );
  ADDFXL mult_241_5_U8 ( .A(mult_241_5_n21), .B(mult_241_5_n22), .CI(
        mult_241_5_n8), .CO(mult_241_5_n7), .S(N1426) );
  ADDFXL mult_241_5_U7 ( .A(mult_241_5_n19), .B(mult_241_5_n20), .CI(
        mult_241_5_n7), .CO(mult_241_5_n6), .S(N1427) );
  ADDFXL mult_241_5_U6 ( .A(mult_241_5_n17), .B(mult_241_5_n18), .CI(
        mult_241_5_n6), .CO(mult_241_5_n5), .S(N1428) );
  ADDFXL mult_241_5_U5 ( .A(mult_241_5_n15), .B(mult_241_5_n16), .CI(
        mult_241_5_n5), .CO(mult_241_5_n4), .S(N1429) );
  ADDFXL mult_241_5_U4 ( .A(mult_241_5_n14), .B(mult_241_5_n13), .CI(
        mult_241_5_n4), .CO(mult_241_5_n3), .S(N1430) );
  ADDFXL mult_241_5_U3 ( .A(mult_241_5_n11), .B(mult_241_5_n12), .CI(
        mult_241_5_n3), .CO(mult_241_5_n2), .S(N1431) );
  ADDFXL mult_241_5_U2 ( .A(mult_241_5_n10), .B(array[157]), .CI(mult_241_5_n2), .CO(N1433), .S(N1432) );
  ADDHXL mult_241_U17 ( .A(array[183]), .B(N13070), .CO(mult_241_n22), .S(
        mult_241_n23) );
  ADDFXL mult_241_U16 ( .A(N13070), .B(array[184]), .CI(array[182]), .CO(
        mult_241_n20), .S(mult_241_n21) );
  ADDFXL mult_241_U15 ( .A(array[182]), .B(array[185]), .CI(array[183]), .CO(
        mult_241_n18), .S(mult_241_n19) );
  ADDFXL mult_241_U14 ( .A(array[183]), .B(array[186]), .CI(array[184]), .CO(
        mult_241_n16), .S(mult_241_n17) );
  ADDFXL mult_241_U13 ( .A(array[184]), .B(array[187]), .CI(array[185]), .CO(
        mult_241_n14), .S(mult_241_n15) );
  ADDHXL mult_241_U12 ( .A(array[186]), .B(array[185]), .CO(mult_241_n12), .S(
        mult_241_n13) );
  ADDHXL mult_241_U11 ( .A(array[187]), .B(array[186]), .CO(mult_241_n10), .S(
        mult_241_n11) );
  ADDHXL mult_241_U10 ( .A(N13060), .B(array[182]), .CO(mult_241_n9), .S(
        N13080) );
  ADDFXL mult_241_U9 ( .A(mult_241_n9), .B(N13060), .CI(mult_241_n23), .CO(
        mult_241_n8), .S(N13090) );
  ADDFXL mult_241_U8 ( .A(mult_241_n21), .B(mult_241_n22), .CI(mult_241_n8), 
        .CO(mult_241_n7), .S(N13100) );
  ADDFXL mult_241_U7 ( .A(mult_241_n19), .B(mult_241_n20), .CI(mult_241_n7), 
        .CO(mult_241_n6), .S(N13110) );
  ADDFXL mult_241_U6 ( .A(mult_241_n17), .B(mult_241_n18), .CI(mult_241_n6), 
        .CO(mult_241_n5), .S(N13120) );
  ADDFXL mult_241_U5 ( .A(mult_241_n15), .B(mult_241_n16), .CI(mult_241_n5), 
        .CO(mult_241_n4), .S(N13130) );
  ADDFXL mult_241_U4 ( .A(mult_241_n14), .B(mult_241_n13), .CI(mult_241_n4), 
        .CO(mult_241_n3), .S(N13140) );
  ADDFXL mult_241_U3 ( .A(mult_241_n11), .B(mult_241_n12), .CI(mult_241_n3), 
        .CO(mult_241_n2), .S(N13150) );
  ADDFXL mult_241_U2 ( .A(mult_241_n10), .B(array[187]), .CI(mult_241_n2), 
        .CO(N13170), .S(N13160) );
  DFFQX1 prev_orig_addr_reg_7_ ( .D(n750), .CK(clk), .Q(n1296) );
  DFFQX1 prev_orig_addr_reg_0_ ( .D(n757), .CK(clk), .Q(N164) );
  DFFQX1 prev_orig_addr_reg_2_ ( .D(n755), .CK(clk), .Q(N668) );
  DFFQX1 i_reg_1_ ( .D(n764), .CK(clk), .Q(i[1]) );
  DFFQX1 i_reg_7_ ( .D(n758), .CK(clk), .Q(i[7]) );
  DFFQX1 i_reg_6_ ( .D(n759), .CK(clk), .Q(i[6]) );
  DFFQX1 i_reg_3_ ( .D(n762), .CK(clk), .Q(i[3]) );
  DFFQX1 i_reg_4_ ( .D(n761), .CK(clk), .Q(i[4]) );
  DFFQX1 i_reg_5_ ( .D(n760), .CK(clk), .Q(i[5]) );
  DFFQX1 j_reg_7_ ( .D(n767), .CK(clk), .Q(j[7]) );
  DFFQX1 j_reg_2_ ( .D(n766), .CK(clk), .Q(j[2]) );
  DFFQX1 j_reg_5_ ( .D(n769), .CK(clk), .Q(j[5]) );
  DFFQX1 j_reg_6_ ( .D(n768), .CK(clk), .Q(j[6]) );
  DFFQX1 j_reg_4_ ( .D(n770), .CK(clk), .Q(j[4]) );
  DFFQX1 j_reg_3_ ( .D(n771), .CK(clk), .Q(j[3]) );
  DFFX1 array_reg_0__1__7_ ( .D(n592), .CK(clk), .Q(array[181]), .QN(n1760) );
  EDFFX1 array_reg_3__4__7_ ( .D(orig_data[7]), .E(n12720), .CK(clk), .Q(
        array[43]), .QN(n320) );
  DFFX1 array_reg_0__1__5_ ( .D(n594), .CK(clk), .Q(array[179]), .QN(n1780) );
  EDFFX1 array_reg_1__4__7_ ( .D(orig_data[7]), .E(n12740), .CK(clk), .Q(
        array[121]), .QN(n240) );
  EDFFX1 array_reg_0__4__7_ ( .D(orig_data[7]), .E(n12750), .CK(clk), .Q(
        array[157]), .QN(n200) );
  DFFX1 array_reg_0__1__6_ ( .D(n593), .CK(clk), .Q(array[180]), .QN(n1770) );
  EDFFX1 array_reg_1__4__6_ ( .D(orig_data[6]), .E(n12740), .CK(clk), .Q(
        array[120]), .QN(n241) );
  EDFFX1 array_reg_3__4__6_ ( .D(orig_data[6]), .E(n12720), .CK(clk), .Q(
        array[42]), .QN(n321) );
  EDFFX1 array_reg_1__4__5_ ( .D(orig_data[5]), .E(n12740), .CK(clk), .Q(
        array[119]), .QN(n242) );
  EDFFX1 array_reg_3__4__5_ ( .D(orig_data[5]), .E(n12720), .CK(clk), .Q(
        array[41]), .QN(n322) );
  DFFX1 array_reg_0__1__4_ ( .D(n595), .CK(clk), .Q(array[178]), .QN(n1790) );
  EDFFX1 array_reg_3__4__4_ ( .D(orig_data[4]), .E(n12720), .CK(clk), .Q(
        array[40]), .QN(n323) );
  DFFX1 array_reg_0__0__7_ ( .D(n584), .CK(clk), .Q(array[187]), .QN(n1680) );
  EDFFX1 array_reg_4__4__7_ ( .D(orig_data[7]), .E(n12710), .CK(clk), .Q(
        array[5]), .QN(n360) );
  DFFX1 array_reg_0__0__6_ ( .D(n585), .CK(clk), .Q(array[186]), .QN(n1690) );
  EDFFX1 array_reg_0__4__6_ ( .D(orig_data[6]), .E(n12750), .CK(clk), .Q(
        array[156]), .QN(n201) );
  EDFFX1 array_reg_4__4__6_ ( .D(orig_data[6]), .E(n12710), .CK(clk), .Q(
        array[4]), .QN(n361) );
  DFFX1 array_reg_0__2__7_ ( .D(n600), .CK(clk), .Q(array[173]), .QN(n1840) );
  DFFX1 array_reg_0__3__3_ ( .D(n612), .CK(clk), .Q(array[161]), .QN(n1960) );
  DFFX1 array_reg_0__1__3_ ( .D(n596), .CK(clk), .Q(array[177]), .QN(n1800) );
  EDFFX1 array_reg_1__4__4_ ( .D(orig_data[4]), .E(n12740), .CK(clk), .Q(
        array[118]), .QN(n243) );
  EDFFX1 array_reg_1__4__3_ ( .D(orig_data[3]), .E(n12740), .CK(clk), .Q(
        array[117]), .QN(n244) );
  EDFFX1 array_reg_3__4__3_ ( .D(orig_data[3]), .E(n12720), .CK(clk), .Q(
        array[39]), .QN(n324) );
  DFFX1 array_reg_0__1__1_ ( .D(n598), .CK(clk), .Q(array[175]), .QN(n1820) );
  DFFX1 array_reg_0__0__5_ ( .D(n586), .CK(clk), .Q(array[185]), .QN(n1700) );
  EDFFX1 array_reg_0__4__5_ ( .D(orig_data[5]), .E(n12750), .CK(clk), .Q(
        array[155]), .QN(n202) );
  EDFFX1 array_reg_4__4__5_ ( .D(orig_data[5]), .E(n12710), .CK(clk), .Q(
        array[3]), .QN(n362) );
  DFFX1 array_reg_0__3__2_ ( .D(n613), .CK(clk), .Q(array[160]), .QN(n1970) );
  DFFX1 array_reg_0__1__2_ ( .D(n597), .CK(clk), .Q(array[176]), .QN(n1810) );
  DFFX1 array_reg_0__1__0_ ( .D(n599), .CK(clk), .Q(array[174]), .QN(n1830) );
  EDFFX1 array_reg_3__4__2_ ( .D(orig_data[2]), .E(n12720), .CK(clk), .Q(
        array[38]), .QN(n325) );
  DFFX1 array_reg_0__2__6_ ( .D(n601), .CK(clk), .Q(array[172]), .QN(n1850) );
  EDFFX1 array_reg_2__4__7_ ( .D(orig_data[7]), .E(n12730), .CK(clk), .Q(
        array[81]), .QN(n280) );
  DFFX1 array_reg_0__3__1_ ( .D(n614), .CK(clk), .Q(array[159]), .QN(n1980) );
  EDFFX1 array_reg_1__4__1_ ( .D(orig_data[1]), .E(n12740), .CK(clk), .Q(
        array[115]), .QN(n246) );
  EDFFX1 array_reg_3__4__1_ ( .D(orig_data[1]), .E(n12720), .CK(clk), .Q(
        array[37]), .QN(n326) );
  DFFX1 array_reg_0__0__4_ ( .D(n587), .CK(clk), .Q(array[184]), .QN(n1710) );
  DFFX1 array_reg_0__0__3_ ( .D(n588), .CK(clk), .Q(array[183]), .QN(n1720) );
  EDFFX1 array_reg_0__4__4_ ( .D(orig_data[4]), .E(n12750), .CK(clk), .Q(
        array[154]), .QN(n203) );
  EDFFX1 array_reg_4__4__4_ ( .D(orig_data[4]), .E(n12710), .CK(clk), .Q(
        array[2]), .QN(n363) );
  EDFFX1 array_reg_0__4__3_ ( .D(orig_data[3]), .E(n12750), .CK(clk), .Q(
        array[153]), .QN(n204) );
  EDFFX1 array_reg_4__4__3_ ( .D(orig_data[3]), .E(n12710), .CK(clk), .Q(
        array[1]), .QN(n364) );
  DFFX1 array_reg_0__0__2_ ( .D(n589), .CK(clk), .Q(array[182]), .QN(n1730) );
  EDFFX1 array_reg_0__4__2_ ( .D(orig_data[2]), .E(n12750), .CK(clk), .Q(
        array[152]), .QN(n205) );
  EDFFX1 array_reg_4__4__2_ ( .D(orig_data[2]), .E(n12710), .CK(clk), .Q(
        array[0]), .QN(n365) );
  DFFX1 array_reg_0__3__0_ ( .D(n615), .CK(clk), .Q(array[158]), .QN(n1990) );
  EDFFX1 array_reg_1__4__2_ ( .D(orig_data[2]), .E(n12740), .CK(clk), .Q(
        array[116]), .QN(n245) );
  EDFFX1 array_reg_1__4__0_ ( .D(orig_data[0]), .E(n12740), .CK(clk), .Q(
        array[114]), .QN(n247) );
  EDFFX1 array_reg_0__4__1_ ( .D(orig_data[1]), .E(n12750), .CK(clk), .Q(N1423), .QN(n206) );
  EDFFX1 array_reg_2__4__6_ ( .D(orig_data[6]), .E(n12730), .CK(clk), .Q(
        array[80]), .QN(n281) );
  DFFX1 array_reg_0__2__4_ ( .D(n603), .CK(clk), .Q(array[170]), .QN(n1870) );
  EDFFX1 array_reg_4__4__0_ ( .D(orig_data[0]), .E(n12710), .CK(clk), .Q(N2226), .QN(n367) );
  DFFX1 array_reg_0__2__5_ ( .D(n602), .CK(clk), .Q(array[171]), .QN(n1860) );
  EDFFX1 array_reg_2__4__5_ ( .D(orig_data[5]), .E(n12730), .CK(clk), .Q(
        array[79]), .QN(n282) );
  DFFX1 array_reg_0__0__1_ ( .D(n590), .CK(clk), .Q(N13070), .QN(n1740) );
  EDFFX1 array_reg_0__4__0_ ( .D(orig_data[0]), .E(n12750), .CK(clk), .Q(N1422), .QN(n207) );
  EDFFX1 array_reg_4__4__1_ ( .D(orig_data[1]), .E(n12710), .CK(clk), .Q(N2227), .QN(n366) );
  EDFFX1 array_reg_3__4__0_ ( .D(orig_data[0]), .E(n12720), .CK(clk), .Q(
        array[36]), .QN(n327) );
  DFFX1 array_reg_0__2__3_ ( .D(n604), .CK(clk), .Q(array[169]), .QN(n1880) );
  EDFFX1 array_reg_2__4__3_ ( .D(orig_data[3]), .E(n12730), .CK(clk), .Q(
        array[77]), .QN(n284) );
  DFFX1 array_reg_0__2__1_ ( .D(n606), .CK(clk), .Q(array[167]), .QN(n1900) );
  EDFFX1 array_reg_2__4__4_ ( .D(orig_data[4]), .E(n12730), .CK(clk), .Q(
        array[78]), .QN(n283) );
  DFFX1 array_reg_0__0__0_ ( .D(n591), .CK(clk), .Q(N13060), .QN(n1750) );
  DFFX1 array_reg_0__2__2_ ( .D(n605), .CK(clk), .Q(array[168]), .QN(n1890) );
  EDFFX1 array_reg_2__4__2_ ( .D(orig_data[2]), .E(n12730), .CK(clk), .Q(
        array[76]), .QN(n285) );
  EDFFX1 array_reg_2__4__1_ ( .D(orig_data[1]), .E(n12730), .CK(clk), .Q(
        array[75]), .QN(n286) );
  EDFFX2 array_reg_2__4__0_ ( .D(orig_data[0]), .E(n12730), .CK(clk), .Q(
        array[74]), .QN(n287) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_14 ( .A(N1332), .B(N2121), .CI(
        add_21_root_add_0_root_add_245_5_carry[14]), .CO(
        add_21_root_add_0_root_add_245_5_carry[15]), .S(N1981) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_14 ( .A(N18800), .B(N1400), .CI(
        add_20_root_add_0_root_add_245_5_carry[14]), .CO(
        add_20_root_add_0_root_add_245_5_carry[15]), .S(N1566) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_15 ( .A(N1881), .B(N1401), .CI(
        add_20_root_add_0_root_add_245_5_carry[15]), .CO(N1568), .S(N1567) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_15 ( .A(N1333), .B(N2122), .CI(
        add_21_root_add_0_root_add_245_5_carry[15]), .CO(N1983), .S(N1982) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_14 ( .A(N2046), .B(N1631), .CI(
        add_18_root_add_0_root_add_245_5_carry[14]), .CO(
        add_18_root_add_0_root_add_245_5_carry[15]), .S(N1938) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_15 ( .A(N2047), .B(N1632), .CI(
        add_18_root_add_0_root_add_245_5_carry[15]), .CO(N19400), .S(N1939) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_14 ( .A(N2200), .B(N1468), .CI(
        add_19_root_add_0_root_add_245_5_carry[14]), .CO(
        add_19_root_add_0_root_add_245_5_carry[15]), .S(N1524) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_15 ( .A(N2201), .B(N1469), .CI(
        add_19_root_add_0_root_add_245_5_carry[15]), .CO(N1526), .S(N1525) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_5 ( .A(
        add_6_root_add_0_root_add_245_5_A_5_), .B(N1744), .CI(
        add_6_root_add_0_root_add_245_5_carry_5_), .CO(
        add_6_root_add_0_root_add_245_5_carry_6_), .S(N1765) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_16 ( .A(N1367), .B(N1672), .CI(
        add_17_root_add_0_root_add_245_5_carry[16]), .CO(N2140), .S(N2139) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_4 ( .A(
        add_6_root_add_0_root_add_245_5_A_4_), .B(N1743), .CI(n807), .CO(
        add_6_root_add_0_root_add_245_5_carry_5_), .S(N1764) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_2 ( .A(N2073), .B(N13070), .CI(
        n803), .CO(add_23_root_add_0_root_add_245_5_carry[3]), .S(N1635) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_2 ( .A(N1423), .B(N2227), .CI(
        n801), .CO(add_22_root_add_0_root_add_245_5_carry[3]), .S(N1596) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_1 ( .A(N1352), .B(N1657), .CI(
        n799), .CO(add_17_root_add_0_root_add_245_5_carry[2]), .S(N1804) );
  DFFQX1 i_reg_2_ ( .D(n763), .CK(clk), .Q(i[2]) );
  DFFQX1 j_reg_1_ ( .D(n772), .CK(clk), .Q(j[1]) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_15 ( .A(N1982), .B(N1567), .CI(
        add_8_root_add_0_root_add_245_5_carry_15_), .CO(
        add_8_root_add_0_root_add_245_5_carry_16_), .S(
        add_6_root_add_0_root_add_245_5_A_15_) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_14 ( .A(N1981), .B(N1566), .CI(
        add_8_root_add_0_root_add_245_5_carry_14_), .CO(
        add_8_root_add_0_root_add_245_5_carry_15_), .S(
        add_6_root_add_0_root_add_245_5_A_14_) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_16 ( .A(N1983), .B(N1568), .CI(
        add_8_root_add_0_root_add_245_5_carry_16_), .CO(
        add_6_root_add_0_root_add_245_5_A_17_), .S(
        add_6_root_add_0_root_add_245_5_A_16_) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_13 ( .A(N1331), .B(N2120), .CI(
        add_21_root_add_0_root_add_245_5_carry[13]), .CO(
        add_21_root_add_0_root_add_245_5_carry[14]), .S(N19800) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_13 ( .A(N1879), .B(N1399), .CI(
        add_20_root_add_0_root_add_245_5_carry[13]), .CO(
        add_20_root_add_0_root_add_245_5_carry[14]), .S(N1565) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_12 ( .A(N1878), .B(N1398), .CI(
        add_20_root_add_0_root_add_245_5_carry[12]), .CO(
        add_20_root_add_0_root_add_245_5_carry[13]), .S(N1564) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_8 ( .A(
        add_6_root_add_0_root_add_245_5_A_8_), .B(N1747), .CI(
        add_6_root_add_0_root_add_245_5_carry_8_), .CO(
        add_6_root_add_0_root_add_245_5_carry_9_), .S(N1768) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_13 ( .A(N2045), .B(N1630), .CI(
        add_18_root_add_0_root_add_245_5_carry[13]), .CO(
        add_18_root_add_0_root_add_245_5_carry[14]), .S(N1937) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_12 ( .A(N2044), .B(N1629), .CI(
        add_18_root_add_0_root_add_245_5_carry[12]), .CO(
        add_18_root_add_0_root_add_245_5_carry[13]), .S(N1936) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_12 ( .A(N1330), .B(N2119), .CI(
        add_21_root_add_0_root_add_245_5_carry[12]), .CO(
        add_21_root_add_0_root_add_245_5_carry[13]), .S(N1979) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_11 ( .A(N2043), .B(N1628), .CI(
        add_18_root_add_0_root_add_245_5_carry[11]), .CO(
        add_18_root_add_0_root_add_245_5_carry[12]), .S(N1935) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_11 ( .A(N1329), .B(N2118), .CI(
        add_21_root_add_0_root_add_245_5_carry[11]), .CO(
        add_21_root_add_0_root_add_245_5_carry[12]), .S(N1978) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_12 ( .A(N2083), .B(N13170), .CI(
        add_23_root_add_0_root_add_245_5_carry[12]), .CO(N1646), .S(N1645) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_13 ( .A(N2199), .B(N1467), .CI(
        add_19_root_add_0_root_add_245_5_carry[13]), .CO(
        add_19_root_add_0_root_add_245_5_carry[14]), .S(N1523) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_12 ( .A(N2198), .B(N1466), .CI(
        add_19_root_add_0_root_add_245_5_carry[12]), .CO(
        add_19_root_add_0_root_add_245_5_carry[13]), .S(N1522) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_11 ( .A(N2197), .B(N1465), .CI(
        add_19_root_add_0_root_add_245_5_carry[11]), .CO(
        add_19_root_add_0_root_add_245_5_carry[12]), .S(N1521) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_11 ( .A(N1877), .B(N1397), .CI(
        add_20_root_add_0_root_add_245_5_carry[11]), .CO(
        add_20_root_add_0_root_add_245_5_carry[12]), .S(N1563) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_12 ( .A(N1433), .B(N2237), .CI(
        add_22_root_add_0_root_add_245_5_carry[12]), .CO(N1607), .S(N1606) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_15 ( .A(N1939), .B(N2138), .CI(
        add_7_root_add_0_root_add_245_5_carry_15_), .CO(
        add_7_root_add_0_root_add_245_5_carry_16_), .S(N1818) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_15 ( .A(N1485), .B(N1525), .CI(
        add_13_root_add_0_root_add_245_5_carry_15_), .CO(
        add_13_root_add_0_root_add_245_5_carry_16_), .S(
        add_13_root_add_0_root_add_245_5_SUM_15_) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_14 ( .A(N1938), .B(N2137), .CI(
        add_7_root_add_0_root_add_245_5_carry_14_), .CO(
        add_7_root_add_0_root_add_245_5_carry_15_), .S(N1817) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_14 ( .A(N1484), .B(N1524), .CI(
        add_13_root_add_0_root_add_245_5_carry_14_), .CO(
        add_13_root_add_0_root_add_245_5_carry_15_), .S(
        add_13_root_add_0_root_add_245_5_SUM_14_) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_7 ( .A(
        add_6_root_add_0_root_add_245_5_A_7_), .B(N1746), .CI(
        add_6_root_add_0_root_add_245_5_carry_7_), .CO(
        add_6_root_add_0_root_add_245_5_carry_8_), .S(N1767) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_6 ( .A(
        add_6_root_add_0_root_add_245_5_A_6_), .B(N1745), .CI(
        add_6_root_add_0_root_add_245_5_carry_6_), .CO(
        add_6_root_add_0_root_add_245_5_carry_7_), .S(N1766) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_11 ( .A(N2082), .B(N13160), .CI(
        add_23_root_add_0_root_add_245_5_carry[11]), .CO(
        add_23_root_add_0_root_add_245_5_carry[12]), .S(N1644) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_5 ( .A(N1323), .B(N2112), .CI(
        add_21_root_add_0_root_add_245_5_carry[5]), .CO(
        add_21_root_add_0_root_add_245_5_carry[6]), .S(N1972) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_11 ( .A(N1432), .B(N2236), .CI(
        add_22_root_add_0_root_add_245_5_carry[11]), .CO(
        add_22_root_add_0_root_add_245_5_carry[12]), .S(N1605) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_5 ( .A(N1871), .B(N1391), .CI(
        add_20_root_add_0_root_add_245_5_carry[5]), .CO(
        add_20_root_add_0_root_add_245_5_carry[6]), .S(N1557) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_16 ( .A(N19400), .B(N2139), .CI(
        add_7_root_add_0_root_add_245_5_carry_16_), .CO(
        add_7_root_add_0_root_add_245_5_carry_17_), .S(N1819) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_16 ( .A(N1486), .B(N1526), .CI(
        add_13_root_add_0_root_add_245_5_carry_16_), .CO(
        add_13_root_add_0_root_add_245_5_carry_17_), .S(
        add_13_root_add_0_root_add_245_5_SUM_16_) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_5 ( .A(N2037), .B(N1622), .CI(
        add_18_root_add_0_root_add_245_5_carry[5]), .CO(
        add_18_root_add_0_root_add_245_5_carry[6]), .S(N1929) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_4 ( .A(N2075), .B(N13090), .CI(
        add_23_root_add_0_root_add_245_5_carry[4]), .CO(
        add_23_root_add_0_root_add_245_5_carry[5]), .S(N1637) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_4 ( .A(N2036), .B(N1621), .CI(
        n805), .CO(add_18_root_add_0_root_add_245_5_carry[5]), .S(N1928) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_4 ( .A(N1322), .B(N2111), .CI(
        n810), .CO(add_21_root_add_0_root_add_245_5_carry[5]), .S(N1971) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_2 ( .A(N1635), .B(N1596), .CI(
        n802), .CO(add_12_root_add_0_root_add_245_5_carry_3_), .S(
        add_9_root_add_0_root_add_245_5_B_2_) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_5 ( .A(N2191), .B(N1459), .CI(
        add_19_root_add_0_root_add_245_5_carry[5]), .CO(
        add_19_root_add_0_root_add_245_5_carry[6]), .S(N1515) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_4 ( .A(N1425), .B(N2229), .CI(
        add_22_root_add_0_root_add_245_5_carry[4]), .CO(
        add_22_root_add_0_root_add_245_5_carry[5]), .S(N1598) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_4 ( .A(N2190), .B(N1458), .CI(
        n804), .CO(add_19_root_add_0_root_add_245_5_carry[5]), .S(N1514) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_4 ( .A(N18700), .B(N1390), .CI(
        n809), .CO(add_20_root_add_0_root_add_245_5_carry[5]), .S(N1556) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_3 ( .A(N1424), .B(N2228), .CI(
        add_22_root_add_0_root_add_245_5_carry[3]), .CO(
        add_22_root_add_0_root_add_245_5_carry[4]), .S(N1597) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_3 ( .A(N2074), .B(N13080), .CI(
        add_23_root_add_0_root_add_245_5_carry[3]), .CO(
        add_23_root_add_0_root_add_245_5_carry[4]), .S(N1636) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_2 ( .A(N1353), .B(N1658), .CI(
        add_17_root_add_0_root_add_245_5_carry[2]), .CO(
        add_17_root_add_0_root_add_245_5_carry[3]), .S(N1805) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_3 ( .A(N1354), .B(N1659), .CI(
        add_17_root_add_0_root_add_245_5_carry[3]), .CO(
        add_17_root_add_0_root_add_245_5_carry[4]), .S(N2126) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_2 ( .A(
        add_9_root_add_0_root_add_245_5_A_2_), .B(
        add_9_root_add_0_root_add_245_5_B_2_), .CI(n800), .CO(
        add_9_root_add_0_root_add_245_5_carry_3_), .S(N2204) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_5 ( .A(N1356), .B(N1661), .CI(
        add_17_root_add_0_root_add_245_5_carry[5]), .CO(
        add_17_root_add_0_root_add_245_5_carry[6]), .S(N2128) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_4 ( .A(N1355), .B(N16600), .CI(
        add_17_root_add_0_root_add_245_5_carry[4]), .CO(
        add_17_root_add_0_root_add_245_5_carry[5]), .S(N2127) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_16 ( .A(
        add_6_root_add_0_root_add_245_5_A_16_), .B(N1755), .CI(
        add_6_root_add_0_root_add_245_5_carry_16_), .CO(
        add_6_root_add_0_root_add_245_5_carry_17_), .S(N1776) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_14 ( .A(
        add_6_root_add_0_root_add_245_5_A_14_), .B(N1753), .CI(
        add_6_root_add_0_root_add_245_5_carry_14_), .CO(
        add_6_root_add_0_root_add_245_5_carry_15_), .S(N1774) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_17 ( .A(
        add_6_root_add_0_root_add_245_5_A_17_), .B(N1756), .CI(
        add_6_root_add_0_root_add_245_5_carry_17_), .CO(
        add_6_root_add_0_root_add_245_5_carry_18_), .S(N1777) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_15 ( .A(
        add_6_root_add_0_root_add_245_5_A_15_), .B(N1754), .CI(
        add_6_root_add_0_root_add_245_5_carry_15_), .CO(
        add_6_root_add_0_root_add_245_5_carry_16_), .S(N1775) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_13 ( .A(
        add_6_root_add_0_root_add_245_5_A_13_), .B(N1752), .CI(
        add_6_root_add_0_root_add_245_5_carry_13_), .CO(
        add_6_root_add_0_root_add_245_5_carry_14_), .S(N1773) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_13 ( .A(N19800), .B(N1565), .CI(
        add_8_root_add_0_root_add_245_5_carry_13_), .CO(
        add_8_root_add_0_root_add_245_5_carry_14_), .S(
        add_6_root_add_0_root_add_245_5_A_13_) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_12 ( .A(
        add_6_root_add_0_root_add_245_5_A_12_), .B(N1751), .CI(
        add_6_root_add_0_root_add_245_5_carry_12_), .CO(
        add_6_root_add_0_root_add_245_5_carry_13_), .S(N1772) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_11 ( .A(
        add_6_root_add_0_root_add_245_5_A_11_), .B(N17500), .CI(
        add_6_root_add_0_root_add_245_5_carry_11_), .CO(
        add_6_root_add_0_root_add_245_5_carry_12_), .S(N1771) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_12 ( .A(N1979), .B(N1564), .CI(
        add_8_root_add_0_root_add_245_5_carry_12_), .CO(
        add_8_root_add_0_root_add_245_5_carry_13_), .S(
        add_6_root_add_0_root_add_245_5_A_12_) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_11 ( .A(N1978), .B(N1563), .CI(
        add_8_root_add_0_root_add_245_5_carry_11_), .CO(
        add_8_root_add_0_root_add_245_5_carry_12_), .S(
        add_6_root_add_0_root_add_245_5_A_11_) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_10 ( .A(
        add_6_root_add_0_root_add_245_5_A_10_), .B(N1749), .CI(
        add_6_root_add_0_root_add_245_5_carry_10_), .CO(
        add_6_root_add_0_root_add_245_5_carry_11_), .S(N17700) );
  ADDFXL add_6_root_add_0_root_add_245_5_U1_9 ( .A(
        add_6_root_add_0_root_add_245_5_A_9_), .B(N1748), .CI(
        add_6_root_add_0_root_add_245_5_carry_9_), .CO(
        add_6_root_add_0_root_add_245_5_carry_10_), .S(N1769) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_10 ( .A(N1328), .B(N2117), .CI(
        add_21_root_add_0_root_add_245_5_carry[10]), .CO(
        add_21_root_add_0_root_add_245_5_carry[11]), .S(N1977) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_9 ( .A(N1327), .B(N2116), .CI(
        add_21_root_add_0_root_add_245_5_carry[9]), .CO(
        add_21_root_add_0_root_add_245_5_carry[10]), .S(N1976) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_8 ( .A(N1326), .B(N2115), .CI(
        add_21_root_add_0_root_add_245_5_carry[8]), .CO(
        add_21_root_add_0_root_add_245_5_carry[9]), .S(N1975) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_13 ( .A(N1646), .B(N1607), .CI(
        add_12_root_add_0_root_add_245_5_carry_13_), .CO(
        add_9_root_add_0_root_add_245_5_B_14_), .S(
        add_9_root_add_0_root_add_245_5_B_13_) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_12 ( .A(N1645), .B(N1606), .CI(
        add_12_root_add_0_root_add_245_5_carry_12_), .CO(
        add_12_root_add_0_root_add_245_5_carry_13_), .S(
        add_9_root_add_0_root_add_245_5_B_12_) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_10 ( .A(N2196), .B(N1464), .CI(
        add_19_root_add_0_root_add_245_5_carry[10]), .CO(
        add_19_root_add_0_root_add_245_5_carry[11]), .S(N1520) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_10 ( .A(N1876), .B(N1396), .CI(
        add_20_root_add_0_root_add_245_5_carry[10]), .CO(
        add_20_root_add_0_root_add_245_5_carry[11]), .S(N1562) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_9 ( .A(N1875), .B(N1395), .CI(
        add_20_root_add_0_root_add_245_5_carry[9]), .CO(
        add_20_root_add_0_root_add_245_5_carry[10]), .S(N1561) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_8 ( .A(N1874), .B(N1394), .CI(
        add_20_root_add_0_root_add_245_5_carry[8]), .CO(
        add_20_root_add_0_root_add_245_5_carry[9]), .S(N1560) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_13 ( .A(N1937), .B(N2136), .CI(
        add_7_root_add_0_root_add_245_5_carry_13_), .CO(
        add_7_root_add_0_root_add_245_5_carry_14_), .S(N1816) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_12 ( .A(N1936), .B(N2135), .CI(
        add_7_root_add_0_root_add_245_5_carry_12_), .CO(
        add_7_root_add_0_root_add_245_5_carry_13_), .S(N1815) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_11 ( .A(N1935), .B(N2134), .CI(
        add_7_root_add_0_root_add_245_5_carry_11_), .CO(
        add_7_root_add_0_root_add_245_5_carry_12_), .S(N1814) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_5 ( .A(N1972), .B(N1557), .CI(
        add_8_root_add_0_root_add_245_5_carry_5_), .CO(
        add_8_root_add_0_root_add_245_5_carry_6_), .S(
        add_6_root_add_0_root_add_245_5_A_5_) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_10 ( .A(N2081), .B(N13150), .CI(
        add_23_root_add_0_root_add_245_5_carry[10]), .CO(
        add_23_root_add_0_root_add_245_5_carry[11]), .S(N1643) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_10 ( .A(N2042), .B(N1627), .CI(
        add_18_root_add_0_root_add_245_5_carry[10]), .CO(
        add_18_root_add_0_root_add_245_5_carry[11]), .S(N1934) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_9 ( .A(N2080), .B(N13140), .CI(
        add_23_root_add_0_root_add_245_5_carry[9]), .CO(
        add_23_root_add_0_root_add_245_5_carry[10]), .S(N1642) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_9 ( .A(N2041), .B(N1626), .CI(
        add_18_root_add_0_root_add_245_5_carry[9]), .CO(
        add_18_root_add_0_root_add_245_5_carry[10]), .S(N1933) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_8 ( .A(N2079), .B(N13130), .CI(
        add_23_root_add_0_root_add_245_5_carry[8]), .CO(
        add_23_root_add_0_root_add_245_5_carry[9]), .S(N1641) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_8 ( .A(N2040), .B(N1625), .CI(
        add_18_root_add_0_root_add_245_5_carry[8]), .CO(
        add_18_root_add_0_root_add_245_5_carry[9]), .S(N1932) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_6 ( .A(N2038), .B(N1623), .CI(
        add_18_root_add_0_root_add_245_5_carry[6]), .CO(
        add_18_root_add_0_root_add_245_5_carry[7]), .S(N19300) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_6 ( .A(N1324), .B(N2113), .CI(
        add_21_root_add_0_root_add_245_5_carry[6]), .CO(
        add_21_root_add_0_root_add_245_5_carry[7]), .S(N1973) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_13 ( .A(
        add_9_root_add_0_root_add_245_5_A_13_), .B(
        add_9_root_add_0_root_add_245_5_B_13_), .CI(
        add_9_root_add_0_root_add_245_5_carry_13_), .CO(
        add_9_root_add_0_root_add_245_5_carry_14_), .S(N2215) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_13 ( .A(N1483), .B(N1523), .CI(
        add_13_root_add_0_root_add_245_5_carry_13_), .CO(
        add_13_root_add_0_root_add_245_5_carry_14_), .S(
        add_13_root_add_0_root_add_245_5_SUM_13_) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_12 ( .A(
        add_9_root_add_0_root_add_245_5_A_12_), .B(
        add_9_root_add_0_root_add_245_5_B_12_), .CI(
        add_9_root_add_0_root_add_245_5_carry_12_), .CO(
        add_9_root_add_0_root_add_245_5_carry_13_), .S(N2214) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_11 ( .A(
        add_9_root_add_0_root_add_245_5_A_11_), .B(
        add_9_root_add_0_root_add_245_5_B_11_), .CI(
        add_9_root_add_0_root_add_245_5_carry_11_), .CO(
        add_9_root_add_0_root_add_245_5_carry_12_), .S(N2213) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_11 ( .A(N1644), .B(N1605), .CI(
        add_12_root_add_0_root_add_245_5_carry_11_), .CO(
        add_12_root_add_0_root_add_245_5_carry_12_), .S(
        add_9_root_add_0_root_add_245_5_B_11_) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_12 ( .A(N1482), .B(N1522), .CI(
        add_13_root_add_0_root_add_245_5_carry_12_), .CO(
        add_13_root_add_0_root_add_245_5_carry_13_), .S(
        add_13_root_add_0_root_add_245_5_SUM_12_) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_11 ( .A(N1481), .B(N1521), .CI(
        add_13_root_add_0_root_add_245_5_carry_11_), .CO(
        add_13_root_add_0_root_add_245_5_carry_12_), .S(
        add_13_root_add_0_root_add_245_5_SUM_11_) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_10 ( .A(
        add_9_root_add_0_root_add_245_5_A_10_), .B(
        add_9_root_add_0_root_add_245_5_B_10_), .CI(
        add_9_root_add_0_root_add_245_5_carry_10_), .CO(
        add_9_root_add_0_root_add_245_5_carry_11_), .S(N2212) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_9 ( .A(
        add_9_root_add_0_root_add_245_5_A_9_), .B(
        add_9_root_add_0_root_add_245_5_B_9_), .CI(
        add_9_root_add_0_root_add_245_5_carry_9_), .CO(
        add_9_root_add_0_root_add_245_5_carry_10_), .S(N2211) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_15 ( .A(N1366), .B(N1671), .CI(
        add_17_root_add_0_root_add_245_5_carry[15]), .CO(
        add_17_root_add_0_root_add_245_5_carry[16]), .S(N2138) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_14 ( .A(N1365), .B(N1670), .CI(
        add_17_root_add_0_root_add_245_5_carry[14]), .CO(
        add_17_root_add_0_root_add_245_5_carry[15]), .S(N2137) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_13 ( .A(N1364), .B(N1669), .CI(
        add_17_root_add_0_root_add_245_5_carry[13]), .CO(
        add_17_root_add_0_root_add_245_5_carry[14]), .S(N2136) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_12 ( .A(N1363), .B(N1668), .CI(
        add_17_root_add_0_root_add_245_5_carry[12]), .CO(
        add_17_root_add_0_root_add_245_5_carry[13]), .S(N2135) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_11 ( .A(N1362), .B(N1667), .CI(
        add_17_root_add_0_root_add_245_5_carry[11]), .CO(
        add_17_root_add_0_root_add_245_5_carry[12]), .S(N2134) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_10 ( .A(N1431), .B(N2235), .CI(
        add_22_root_add_0_root_add_245_5_carry[10]), .CO(
        add_22_root_add_0_root_add_245_5_carry[11]), .S(N1604) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_10 ( .A(N1361), .B(N1666), .CI(
        add_17_root_add_0_root_add_245_5_carry[10]), .CO(
        add_17_root_add_0_root_add_245_5_carry[11]), .S(N2133) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_9 ( .A(N1430), .B(N2234), .CI(
        add_22_root_add_0_root_add_245_5_carry[9]), .CO(
        add_22_root_add_0_root_add_245_5_carry[10]), .S(N1603) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_9 ( .A(N2195), .B(N1463), .CI(
        add_19_root_add_0_root_add_245_5_carry[9]), .CO(
        add_19_root_add_0_root_add_245_5_carry[10]), .S(N1519) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_8 ( .A(N1429), .B(N2233), .CI(
        add_22_root_add_0_root_add_245_5_carry[8]), .CO(
        add_22_root_add_0_root_add_245_5_carry[9]), .S(N1602) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_8 ( .A(N2194), .B(N1462), .CI(
        add_19_root_add_0_root_add_245_5_carry[8]), .CO(
        add_19_root_add_0_root_add_245_5_carry[9]), .S(N1518) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_6 ( .A(N2192), .B(N1460), .CI(
        add_19_root_add_0_root_add_245_5_carry[6]), .CO(
        add_19_root_add_0_root_add_245_5_carry[7]), .S(N1516) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_6 ( .A(N1872), .B(N1392), .CI(
        add_20_root_add_0_root_add_245_5_carry[6]), .CO(
        add_20_root_add_0_root_add_245_5_carry[7]), .S(N1558) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_14 ( .A(
        add_9_root_add_0_root_add_245_5_A_14_), .B(
        add_9_root_add_0_root_add_245_5_B_14_), .CI(
        add_9_root_add_0_root_add_245_5_carry_14_), .CO(
        add_9_root_add_0_root_add_245_5_carry_15_), .S(N2216) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_4 ( .A(N1971), .B(N1556), .CI(n808), .CO(add_8_root_add_0_root_add_245_5_carry_5_), .S(
        add_6_root_add_0_root_add_245_5_A_4_) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_7 ( .A(N2078), .B(N13120), .CI(
        add_23_root_add_0_root_add_245_5_carry[7]), .CO(
        add_23_root_add_0_root_add_245_5_carry[8]), .S(N16400) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_6 ( .A(N2077), .B(N13110), .CI(
        add_23_root_add_0_root_add_245_5_carry[6]), .CO(
        add_23_root_add_0_root_add_245_5_carry[7]), .S(N1639) );
  ADDFXL add_23_root_add_0_root_add_245_5_U1_5 ( .A(N2076), .B(N13100), .CI(
        add_23_root_add_0_root_add_245_5_carry[5]), .CO(
        add_23_root_add_0_root_add_245_5_carry[6]), .S(N1638) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_8 ( .A(
        add_9_root_add_0_root_add_245_5_A_8_), .B(
        add_9_root_add_0_root_add_245_5_B_8_), .CI(
        add_9_root_add_0_root_add_245_5_carry_8_), .CO(
        add_9_root_add_0_root_add_245_5_carry_9_), .S(N2210) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_7 ( .A(
        add_9_root_add_0_root_add_245_5_A_7_), .B(
        add_9_root_add_0_root_add_245_5_B_7_), .CI(
        add_9_root_add_0_root_add_245_5_carry_7_), .CO(
        add_9_root_add_0_root_add_245_5_carry_8_), .S(N2209) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_6 ( .A(
        add_9_root_add_0_root_add_245_5_A_6_), .B(
        add_9_root_add_0_root_add_245_5_B_6_), .CI(
        add_9_root_add_0_root_add_245_5_carry_6_), .CO(
        add_9_root_add_0_root_add_245_5_carry_7_), .S(N2208) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_5 ( .A(
        add_9_root_add_0_root_add_245_5_A_5_), .B(
        add_9_root_add_0_root_add_245_5_B_5_), .CI(
        add_9_root_add_0_root_add_245_5_carry_5_), .CO(
        add_9_root_add_0_root_add_245_5_carry_6_), .S(N2207) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_4 ( .A(N1637), .B(N1598), .CI(
        add_12_root_add_0_root_add_245_5_carry_4_), .CO(
        add_12_root_add_0_root_add_245_5_carry_5_), .S(
        add_9_root_add_0_root_add_245_5_B_4_) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_9 ( .A(N1360), .B(N1665), .CI(
        add_17_root_add_0_root_add_245_5_carry[9]), .CO(
        add_17_root_add_0_root_add_245_5_carry[10]), .S(N2132) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_8 ( .A(N1359), .B(N1664), .CI(
        add_17_root_add_0_root_add_245_5_carry[8]), .CO(
        add_17_root_add_0_root_add_245_5_carry[9]), .S(N2131) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_7 ( .A(N1428), .B(N2232), .CI(
        add_22_root_add_0_root_add_245_5_carry[7]), .CO(
        add_22_root_add_0_root_add_245_5_carry[8]), .S(N1601) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_7 ( .A(N1358), .B(N1663), .CI(
        add_17_root_add_0_root_add_245_5_carry[7]), .CO(
        add_17_root_add_0_root_add_245_5_carry[8]), .S(N2130) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_6 ( .A(N1427), .B(N2231), .CI(
        add_22_root_add_0_root_add_245_5_carry[6]), .CO(
        add_22_root_add_0_root_add_245_5_carry[7]), .S(N1600) );
  ADDFXL add_17_root_add_0_root_add_245_5_U1_6 ( .A(N1357), .B(N1662), .CI(
        add_17_root_add_0_root_add_245_5_carry[6]), .CO(
        add_17_root_add_0_root_add_245_5_carry[7]), .S(N2129) );
  ADDFXL add_22_root_add_0_root_add_245_5_U1_5 ( .A(N1426), .B(N2230), .CI(
        add_22_root_add_0_root_add_245_5_carry[5]), .CO(
        add_22_root_add_0_root_add_245_5_carry[6]), .S(N1599) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_5 ( .A(N1929), .B(N2128), .CI(
        add_7_root_add_0_root_add_245_5_carry_5_), .CO(
        add_7_root_add_0_root_add_245_5_carry_6_), .S(N1808) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_4 ( .A(N1928), .B(N2127), .CI(n798), .CO(add_7_root_add_0_root_add_245_5_carry_5_), .S(N1807) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_5 ( .A(N1475), .B(N1515), .CI(
        add_13_root_add_0_root_add_245_5_carry_5_), .CO(
        add_13_root_add_0_root_add_245_5_carry_6_), .S(
        add_13_root_add_0_root_add_245_5_SUM_5_) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_4 ( .A(
        add_9_root_add_0_root_add_245_5_A_4_), .B(
        add_9_root_add_0_root_add_245_5_B_4_), .CI(
        add_9_root_add_0_root_add_245_5_carry_4_), .CO(
        add_9_root_add_0_root_add_245_5_carry_5_), .S(N2206) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_4 ( .A(N1474), .B(N1514), .CI(
        n797), .CO(add_13_root_add_0_root_add_245_5_carry_5_), .S(
        add_13_root_add_0_root_add_245_5_SUM_4_) );
  ADDFXL add_9_root_add_0_root_add_245_5_U1_3 ( .A(
        add_9_root_add_0_root_add_245_5_A_3_), .B(
        add_9_root_add_0_root_add_245_5_B_3_), .CI(
        add_9_root_add_0_root_add_245_5_carry_3_), .CO(
        add_9_root_add_0_root_add_245_5_carry_4_), .S(N2205) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_3 ( .A(N1636), .B(N1597), .CI(
        add_12_root_add_0_root_add_245_5_carry_3_), .CO(
        add_12_root_add_0_root_add_245_5_carry_4_), .S(
        add_9_root_add_0_root_add_245_5_B_3_) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_10 ( .A(N1977), .B(N1562), .CI(
        add_8_root_add_0_root_add_245_5_carry_10_), .CO(
        add_8_root_add_0_root_add_245_5_carry_11_), .S(
        add_6_root_add_0_root_add_245_5_A_10_) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_9 ( .A(N1976), .B(N1561), .CI(
        add_8_root_add_0_root_add_245_5_carry_9_), .CO(
        add_8_root_add_0_root_add_245_5_carry_10_), .S(
        add_6_root_add_0_root_add_245_5_A_9_) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_8 ( .A(N1975), .B(N1560), .CI(
        add_8_root_add_0_root_add_245_5_carry_8_), .CO(
        add_8_root_add_0_root_add_245_5_carry_9_), .S(
        add_6_root_add_0_root_add_245_5_A_8_) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_10 ( .A(N1934), .B(N2133), .CI(
        add_7_root_add_0_root_add_245_5_carry_10_), .CO(
        add_7_root_add_0_root_add_245_5_carry_11_), .S(N1813) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_6 ( .A(N1973), .B(N1558), .CI(
        add_8_root_add_0_root_add_245_5_carry_6_), .CO(
        add_8_root_add_0_root_add_245_5_carry_7_), .S(
        add_6_root_add_0_root_add_245_5_A_6_) );
  ADDFXL add_18_root_add_0_root_add_245_5_U1_7 ( .A(N2039), .B(N1624), .CI(
        add_18_root_add_0_root_add_245_5_carry[7]), .CO(
        add_18_root_add_0_root_add_245_5_carry[8]), .S(N1931) );
  ADDFXL add_21_root_add_0_root_add_245_5_U1_7 ( .A(N1325), .B(N2114), .CI(
        add_21_root_add_0_root_add_245_5_carry[7]), .CO(
        add_21_root_add_0_root_add_245_5_carry[8]), .S(N1974) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_10 ( .A(N1643), .B(N1604), .CI(
        add_12_root_add_0_root_add_245_5_carry_10_), .CO(
        add_12_root_add_0_root_add_245_5_carry_11_), .S(
        add_9_root_add_0_root_add_245_5_B_10_) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_9 ( .A(N1642), .B(N1603), .CI(
        add_12_root_add_0_root_add_245_5_carry_9_), .CO(
        add_12_root_add_0_root_add_245_5_carry_10_), .S(
        add_9_root_add_0_root_add_245_5_B_9_) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_8 ( .A(N1641), .B(N1602), .CI(
        add_12_root_add_0_root_add_245_5_carry_8_), .CO(
        add_12_root_add_0_root_add_245_5_carry_9_), .S(
        add_9_root_add_0_root_add_245_5_B_8_) );
  ADDFXL add_19_root_add_0_root_add_245_5_U1_7 ( .A(N2193), .B(N1461), .CI(
        add_19_root_add_0_root_add_245_5_carry[7]), .CO(
        add_19_root_add_0_root_add_245_5_carry[8]), .S(N1517) );
  ADDFXL add_20_root_add_0_root_add_245_5_U1_7 ( .A(N1873), .B(N1393), .CI(
        add_20_root_add_0_root_add_245_5_carry[7]), .CO(
        add_20_root_add_0_root_add_245_5_carry[8]), .S(N1559) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_9 ( .A(N1933), .B(N2132), .CI(
        add_7_root_add_0_root_add_245_5_carry_9_), .CO(
        add_7_root_add_0_root_add_245_5_carry_10_), .S(N1812) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_8 ( .A(N1932), .B(N2131), .CI(
        add_7_root_add_0_root_add_245_5_carry_8_), .CO(
        add_7_root_add_0_root_add_245_5_carry_9_), .S(N1811) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_7 ( .A(N1931), .B(N2130), .CI(
        add_7_root_add_0_root_add_245_5_carry_7_), .CO(
        add_7_root_add_0_root_add_245_5_carry_8_), .S(N18100) );
  ADDFXL add_7_root_add_0_root_add_245_5_U1_6 ( .A(N19300), .B(N2129), .CI(
        add_7_root_add_0_root_add_245_5_carry_6_), .CO(
        add_7_root_add_0_root_add_245_5_carry_7_), .S(N1809) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_10 ( .A(N1480), .B(N1520), .CI(
        add_13_root_add_0_root_add_245_5_carry_10_), .CO(
        add_13_root_add_0_root_add_245_5_carry_11_), .S(
        add_13_root_add_0_root_add_245_5_SUM_10_) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_9 ( .A(N1479), .B(N1519), .CI(
        add_13_root_add_0_root_add_245_5_carry_9_), .CO(
        add_13_root_add_0_root_add_245_5_carry_10_), .S(
        add_13_root_add_0_root_add_245_5_SUM_9_) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_8 ( .A(N1478), .B(N1518), .CI(
        add_13_root_add_0_root_add_245_5_carry_8_), .CO(
        add_13_root_add_0_root_add_245_5_carry_9_), .S(
        add_13_root_add_0_root_add_245_5_SUM_8_) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_7 ( .A(N16400), .B(N1601), .CI(
        add_12_root_add_0_root_add_245_5_carry_7_), .CO(
        add_12_root_add_0_root_add_245_5_carry_8_), .S(
        add_9_root_add_0_root_add_245_5_B_7_) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_7 ( .A(N1477), .B(N1517), .CI(
        add_13_root_add_0_root_add_245_5_carry_7_), .CO(
        add_13_root_add_0_root_add_245_5_carry_8_), .S(
        add_13_root_add_0_root_add_245_5_SUM_7_) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_6 ( .A(N1639), .B(N1600), .CI(
        add_12_root_add_0_root_add_245_5_carry_6_), .CO(
        add_12_root_add_0_root_add_245_5_carry_7_), .S(
        add_9_root_add_0_root_add_245_5_B_6_) );
  ADDFXL add_12_root_add_0_root_add_245_5_U1_5 ( .A(N1638), .B(N1599), .CI(
        add_12_root_add_0_root_add_245_5_carry_5_), .CO(
        add_12_root_add_0_root_add_245_5_carry_6_), .S(
        add_9_root_add_0_root_add_245_5_B_5_) );
  ADDFXL add_13_root_add_0_root_add_245_5_U1_6 ( .A(N1476), .B(N1516), .CI(
        add_13_root_add_0_root_add_245_5_carry_6_), .CO(
        add_13_root_add_0_root_add_245_5_carry_7_), .S(
        add_13_root_add_0_root_add_245_5_SUM_6_) );
  ADDFXL add_8_root_add_0_root_add_245_5_U1_7 ( .A(N1974), .B(N1559), .CI(
        add_8_root_add_0_root_add_245_5_carry_7_), .CO(
        add_8_root_add_0_root_add_245_5_carry_8_), .S(
        add_6_root_add_0_root_add_245_5_A_7_) );
  DFFRX1 imgproc_ready_reg ( .D(next_imgproc_ready), .CK(clk), .RN(n971), .QN(
        n795) );
  DFFRX1 request_reg ( .D(next_request), .CK(clk), .RN(n971), .QN(n796) );
  DFFRHQX1 finish_reg ( .D(next_finish), .CK(clk), .RN(n12700), .Q(n848) );
  DFFRX1 row_reg_6_ ( .D(n783), .CK(clk), .RN(n12700), .Q(row[6]), .QN(n1058)
         );
  DFFRX1 row_reg_3_ ( .D(n786), .CK(clk), .RN(n12700), .Q(row[3]), .QN(n1055)
         );
  DFFRX1 row_reg_0_ ( .D(n789), .CK(clk), .RN(n12700), .Q(row[0]), .QN(n1051)
         );
  DFFRX1 row_reg_4_ ( .D(n785), .CK(clk), .RN(n12700), .Q(row[4]), .QN(n1056)
         );
  DFFRX1 row_reg_1_ ( .D(n788), .CK(clk), .RN(n12700), .Q(row[1]), .QN(n1053)
         );
  DFFRX1 row_reg_2_ ( .D(n787), .CK(clk), .RN(n12700), .Q(row[2]), .QN(n1054)
         );
  DFFRX1 row_reg_5_ ( .D(n784), .CK(clk), .RN(n12700), .Q(row[5]), .QN(n1057)
         );
  DFFRX1 row_reg_7_ ( .D(n782), .CK(clk), .RN(n12700), .Q(row[7]), .QN(n1059)
         );
  DFFRX1 state_reg_1_ ( .D(n790), .CK(clk), .RN(n12700), .Q(state[1]), .QN(
        n1065) );
  DFFRX1 state_reg_0_ ( .D(n791), .CK(clk), .RN(n12700), .Q(state[0]) );
  DFFX1 j_reg_0_ ( .D(n773), .CK(clk), .Q(j[0]), .QN(n1218) );
  DFFX1 i_reg_0_ ( .D(n765), .CK(clk), .Q(i[0]), .QN(n1183) );
  DFFX1 array_reg_2__2__5_ ( .D(n666), .CK(clk), .Q(array[95]), .QN(n266) );
  DFFX1 array_reg_2__2__0_ ( .D(n6710), .CK(clk), .Q(array[90]), .QN(n271) );
  DFFX1 array_reg_4__2__7_ ( .D(n728), .CK(clk), .Q(array[21]), .QN(n344) );
  DFFX1 array_reg_4__2__6_ ( .D(n729), .CK(clk), .Q(array[20]), .QN(n345) );
  DFFX1 array_reg_4__2__5_ ( .D(n730), .CK(clk), .Q(array[19]), .QN(n346) );
  DFFX1 array_reg_4__2__4_ ( .D(n731), .CK(clk), .Q(array[18]), .QN(n347) );
  DFFX1 array_reg_4__2__3_ ( .D(n732), .CK(clk), .Q(array[17]), .QN(n348) );
  DFFX1 array_reg_4__2__2_ ( .D(n733), .CK(clk), .Q(array[16]), .QN(n349) );
  DFFX1 array_reg_4__2__1_ ( .D(n734), .CK(clk), .Q(array[15]), .QN(n350) );
  DFFX1 array_reg_4__1__7_ ( .D(n720), .CK(clk), .Q(array[29]), .QN(n336) );
  DFFX1 array_reg_4__1__6_ ( .D(n721), .CK(clk), .Q(array[28]), .QN(n337) );
  DFFX1 array_reg_4__1__5_ ( .D(n722), .CK(clk), .Q(array[27]), .QN(n338) );
  DFFX1 array_reg_4__1__4_ ( .D(n723), .CK(clk), .Q(array[26]), .QN(n339) );
  DFFX1 array_reg_4__1__3_ ( .D(n724), .CK(clk), .Q(array[25]), .QN(n340) );
  DFFX1 array_reg_4__1__2_ ( .D(n725), .CK(clk), .Q(array[24]), .QN(n341) );
  DFFX1 array_reg_4__1__1_ ( .D(n726), .CK(clk), .Q(array[23]), .QN(n342) );
  DFFX1 array_reg_4__1__0_ ( .D(n727), .CK(clk), .Q(array[22]), .QN(n343) );
  DFFX1 array_reg_4__0__7_ ( .D(n712), .CK(clk), .Q(array[35]), .QN(n328) );
  DFFX1 array_reg_4__0__6_ ( .D(n713), .CK(clk), .Q(array[34]), .QN(n329) );
  DFFX1 array_reg_4__0__5_ ( .D(n714), .CK(clk), .Q(array[33]), .QN(n330) );
  DFFX1 array_reg_4__0__4_ ( .D(n715), .CK(clk), .Q(array[32]), .QN(n331) );
  DFFX1 array_reg_4__0__3_ ( .D(n716), .CK(clk), .Q(array[31]), .QN(n332) );
  DFFX1 array_reg_4__0__2_ ( .D(n717), .CK(clk), .Q(array[30]), .QN(n333) );
  DFFX1 array_reg_4__0__1_ ( .D(n718), .CK(clk), .Q(N2073), .QN(n334) );
  DFFX1 array_reg_4__0__0_ ( .D(n719), .CK(clk), .Q(N2072), .QN(n335) );
  DFFX1 array_reg_3__3__7_ ( .D(n704), .CK(clk), .Q(array[50]), .QN(n1011) );
  DFFX1 array_reg_3__3__6_ ( .D(n705), .CK(clk), .Q(array[49]), .QN(n1010) );
  DFFX1 array_reg_3__3__5_ ( .D(n706), .CK(clk), .Q(array[48]), .QN(n1009) );
  DFFX1 array_reg_3__3__4_ ( .D(n707), .CK(clk), .Q(array[47]), .QN(n10080) );
  DFFX1 array_reg_3__3__3_ ( .D(n708), .CK(clk), .Q(array[46]), .QN(n10070) );
  DFFX1 array_reg_3__3__2_ ( .D(n709), .CK(clk), .Q(array[45]), .QN(n10060) );
  DFFX1 array_reg_3__3__1_ ( .D(n710), .CK(clk), .Q(array[44]), .QN(n10050) );
  DFFX1 array_reg_3__3__0_ ( .D(n711), .CK(clk), .Q(N19900), .QN(n10040) );
  DFFX1 array_reg_3__2__7_ ( .D(n696), .CK(clk), .Q(array[58]), .QN(n304) );
  DFFX1 array_reg_3__2__6_ ( .D(n697), .CK(clk), .Q(array[57]), .QN(n305) );
  DFFX1 array_reg_3__2__5_ ( .D(n698), .CK(clk), .Q(array[56]), .QN(n306) );
  DFFX1 array_reg_3__2__4_ ( .D(n699), .CK(clk), .Q(array[55]), .QN(n307) );
  DFFX1 array_reg_3__2__3_ ( .D(n700), .CK(clk), .Q(array[54]), .QN(n308) );
  DFFX1 array_reg_3__2__2_ ( .D(n701), .CK(clk), .Q(array[53]), .QN(n309) );
  DFFX1 array_reg_3__2__1_ ( .D(n702), .CK(clk), .Q(array[52]), .QN(n310) );
  DFFX1 array_reg_3__2__0_ ( .D(n703), .CK(clk), .Q(array[51]), .QN(n311) );
  DFFX1 array_reg_3__1__7_ ( .D(n688), .CK(clk), .Q(array[65]), .QN(n10010) );
  DFFX1 array_reg_3__1__6_ ( .D(n689), .CK(clk), .Q(array[64]), .QN(n10000) );
  DFFX1 array_reg_3__1__5_ ( .D(n690), .CK(clk), .Q(array[63]), .QN(n9990) );
  DFFX1 array_reg_3__1__4_ ( .D(n691), .CK(clk), .Q(array[62]), .QN(n9980) );
  DFFX1 array_reg_3__1__3_ ( .D(n692), .CK(clk), .Q(array[61]), .QN(n9970) );
  DFFX1 array_reg_3__1__2_ ( .D(n693), .CK(clk), .Q(array[60]), .QN(n9960) );
  DFFX1 array_reg_3__1__1_ ( .D(n694), .CK(clk), .Q(array[59]), .QN(n995) );
  DFFX1 array_reg_3__1__0_ ( .D(n695), .CK(clk), .Q(N1905), .QN(n994) );
  DFFX1 array_reg_3__0__7_ ( .D(n680), .CK(clk), .Q(array[73]), .QN(n288) );
  DFFX1 array_reg_3__0__6_ ( .D(n681), .CK(clk), .Q(array[72]), .QN(n289) );
  DFFX1 array_reg_3__0__5_ ( .D(n682), .CK(clk), .Q(array[71]), .QN(n290) );
  DFFX1 array_reg_3__0__4_ ( .D(n683), .CK(clk), .Q(array[70]), .QN(n291) );
  DFFX1 array_reg_3__0__3_ ( .D(n684), .CK(clk), .Q(array[69]), .QN(n292) );
  DFFX1 array_reg_3__0__2_ ( .D(n685), .CK(clk), .Q(array[68]), .QN(n293) );
  DFFX1 array_reg_3__0__1_ ( .D(n686), .CK(clk), .Q(array[67]), .QN(n294) );
  DFFX1 array_reg_3__0__0_ ( .D(n687), .CK(clk), .Q(array[66]), .QN(n295) );
  DFFX1 array_reg_2__2__7_ ( .D(n664), .CK(clk), .Q(array[97]), .QN(n264) );
  DFFX1 array_reg_2__2__6_ ( .D(n665), .CK(clk), .Q(array[96]), .QN(n265) );
  DFFX1 array_reg_2__2__4_ ( .D(n667), .CK(clk), .Q(array[94]), .QN(n267) );
  DFFX1 array_reg_2__2__3_ ( .D(n6680), .CK(clk), .Q(array[93]), .QN(n268) );
  DFFX1 array_reg_2__2__2_ ( .D(n6690), .CK(clk), .Q(array[92]), .QN(n269) );
  DFFX1 array_reg_2__2__1_ ( .D(n6700), .CK(clk), .Q(array[91]), .QN(n270) );
  DFFX1 array_reg_2__1__7_ ( .D(n656), .CK(clk), .Q(array[105]), .QN(n256) );
  DFFX1 array_reg_2__1__6_ ( .D(n657), .CK(clk), .Q(array[104]), .QN(n257) );
  DFFX1 array_reg_2__1__5_ ( .D(n658), .CK(clk), .Q(array[103]), .QN(n258) );
  DFFX1 array_reg_2__1__4_ ( .D(n659), .CK(clk), .Q(array[102]), .QN(n259) );
  DFFX1 array_reg_2__1__3_ ( .D(n660), .CK(clk), .Q(array[101]), .QN(n260) );
  DFFX1 array_reg_2__1__2_ ( .D(n661), .CK(clk), .Q(array[100]), .QN(n261) );
  DFFX1 array_reg_2__1__1_ ( .D(n662), .CK(clk), .Q(array[99]), .QN(n262) );
  DFFX1 array_reg_2__1__0_ ( .D(n663), .CK(clk), .Q(array[98]), .QN(n263) );
  DFFX1 array_reg_2__0__7_ ( .D(n648), .CK(clk), .Q(array[113]), .QN(n248) );
  DFFX1 array_reg_2__0__6_ ( .D(n649), .CK(clk), .Q(array[112]), .QN(n249) );
  DFFX1 array_reg_2__0__5_ ( .D(n650), .CK(clk), .Q(array[111]), .QN(n250) );
  DFFX1 array_reg_2__0__4_ ( .D(n651), .CK(clk), .Q(array[110]), .QN(n251) );
  DFFX1 array_reg_2__0__3_ ( .D(n652), .CK(clk), .Q(array[109]), .QN(n252) );
  DFFX1 array_reg_2__0__2_ ( .D(n653), .CK(clk), .Q(array[108]), .QN(n253) );
  DFFX1 array_reg_2__0__1_ ( .D(n654), .CK(clk), .Q(array[107]), .QN(n254) );
  DFFX1 array_reg_4__3__7_ ( .D(n736), .CK(clk), .Q(array[13]), .QN(n352) );
  DFFX1 array_reg_4__3__6_ ( .D(n737), .CK(clk), .Q(array[12]), .QN(n353) );
  DFFX1 array_reg_4__3__5_ ( .D(n738), .CK(clk), .Q(array[11]), .QN(n354) );
  DFFX1 array_reg_4__3__4_ ( .D(n739), .CK(clk), .Q(array[10]), .QN(n355) );
  DFFX1 array_reg_4__3__3_ ( .D(n740), .CK(clk), .Q(array[9]), .QN(n356) );
  DFFX1 array_reg_4__3__2_ ( .D(n741), .CK(clk), .Q(array[8]), .QN(n357) );
  DFFX1 array_reg_4__3__1_ ( .D(n742), .CK(clk), .Q(array[7]), .QN(n358) );
  DFFX1 array_reg_4__3__0_ ( .D(n743), .CK(clk), .Q(array[6]), .QN(n359) );
  DFFX1 array_reg_2__3__7_ ( .D(n6720), .CK(clk), .Q(array[89]), .QN(n272) );
  DFFX1 array_reg_2__3__6_ ( .D(n6730), .CK(clk), .Q(array[88]), .QN(n273) );
  DFFX1 array_reg_2__3__5_ ( .D(n6740), .CK(clk), .Q(array[87]), .QN(n274) );
  DFFX1 array_reg_2__3__4_ ( .D(n6750), .CK(clk), .Q(array[86]), .QN(n275) );
  DFFX1 array_reg_2__3__3_ ( .D(n6760), .CK(clk), .Q(array[85]), .QN(n276) );
  DFFX1 array_reg_2__3__2_ ( .D(n6770), .CK(clk), .Q(array[84]), .QN(n277) );
  DFFX1 array_reg_2__3__1_ ( .D(n6780), .CK(clk), .Q(array[83]), .QN(n278) );
  DFFX1 array_reg_2__3__0_ ( .D(n6790), .CK(clk), .Q(array[82]), .QN(n279) );
  DFFX1 array_reg_1__3__7_ ( .D(n640), .CK(clk), .Q(array[128]), .QN(n991) );
  DFFX1 array_reg_1__3__6_ ( .D(n641), .CK(clk), .Q(array[127]), .QN(n990) );
  DFFX1 array_reg_1__3__5_ ( .D(n642), .CK(clk), .Q(array[126]), .QN(n989) );
  DFFX1 array_reg_1__3__4_ ( .D(n643), .CK(clk), .Q(array[125]), .QN(n988) );
  DFFX1 array_reg_1__3__3_ ( .D(n644), .CK(clk), .Q(array[124]), .QN(n987) );
  DFFX1 array_reg_1__3__2_ ( .D(n645), .CK(clk), .Q(array[123]), .QN(n986) );
  DFFX1 array_reg_1__3__1_ ( .D(n646), .CK(clk), .Q(array[122]), .QN(n985) );
  DFFX1 array_reg_1__3__0_ ( .D(n647), .CK(clk), .Q(N1575), .QN(n984) );
  DFFX1 array_reg_1__2__7_ ( .D(n632), .CK(clk), .Q(array[136]), .QN(n224) );
  DFFX1 array_reg_1__2__6_ ( .D(n633), .CK(clk), .Q(array[135]), .QN(n225) );
  DFFX1 array_reg_1__2__5_ ( .D(n634), .CK(clk), .Q(array[134]), .QN(n226) );
  DFFX1 array_reg_1__2__4_ ( .D(n635), .CK(clk), .Q(array[133]), .QN(n227) );
  DFFX1 array_reg_1__2__3_ ( .D(n636), .CK(clk), .Q(array[132]), .QN(n228) );
  DFFX1 array_reg_1__2__2_ ( .D(n637), .CK(clk), .Q(array[131]), .QN(n229) );
  DFFX1 array_reg_1__2__1_ ( .D(n638), .CK(clk), .Q(array[130]), .QN(n230) );
  DFFX1 array_reg_1__2__0_ ( .D(n639), .CK(clk), .Q(array[129]), .QN(n231) );
  DFFX1 array_reg_1__1__7_ ( .D(n624), .CK(clk), .Q(array[143]), .QN(n981) );
  DFFX1 array_reg_1__1__6_ ( .D(n625), .CK(clk), .Q(array[142]), .QN(n980) );
  DFFX1 array_reg_1__1__5_ ( .D(n626), .CK(clk), .Q(array[141]), .QN(n979) );
  DFFX1 array_reg_1__1__4_ ( .D(n627), .CK(clk), .Q(array[140]), .QN(n978) );
  DFFX1 array_reg_1__1__3_ ( .D(n628), .CK(clk), .Q(array[139]), .QN(n977) );
  DFFX1 array_reg_1__1__2_ ( .D(n629), .CK(clk), .Q(array[138]), .QN(n976) );
  DFFX1 array_reg_1__1__1_ ( .D(n630), .CK(clk), .Q(array[137]), .QN(n975) );
  DFFX1 array_reg_1__1__0_ ( .D(n631), .CK(clk), .Q(N1491), .QN(n974) );
  DFFX1 array_reg_1__0__7_ ( .D(n616), .CK(clk), .Q(array[151]), .QN(n208) );
  DFFX1 array_reg_1__0__6_ ( .D(n617), .CK(clk), .Q(array[150]), .QN(n209) );
  DFFX1 array_reg_1__0__5_ ( .D(n618), .CK(clk), .Q(array[149]), .QN(n210) );
  DFFX1 array_reg_1__0__4_ ( .D(n619), .CK(clk), .Q(array[148]), .QN(n211) );
  DFFX1 array_reg_1__0__3_ ( .D(n620), .CK(clk), .Q(array[147]), .QN(n212) );
  DFFX1 array_reg_1__0__2_ ( .D(n621), .CK(clk), .Q(array[146]), .QN(n213) );
  DFFX1 array_reg_1__0__1_ ( .D(n622), .CK(clk), .Q(array[145]), .QN(n214) );
  DFFX1 array_reg_1__0__0_ ( .D(n623), .CK(clk), .Q(array[144]), .QN(n215) );
  DFFX1 array_reg_0__3__7_ ( .D(n608), .CK(clk), .Q(array[165]), .QN(n1920) );
  DFFX1 array_reg_0__3__6_ ( .D(n609), .CK(clk), .Q(array[164]), .QN(n1930) );
  DFFX1 array_reg_0__3__5_ ( .D(n610), .CK(clk), .Q(array[163]), .QN(n1940) );
  DFFX1 array_reg_0__3__4_ ( .D(n611), .CK(clk), .Q(array[162]), .QN(n1950) );
  DFFSRXL imgproc_addr_reg_6_ ( .D(n576), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1304), .QN(n1241) );
  DFFSRXL imgproc_addr_reg_5_ ( .D(n575), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1305), .QN(n1240) );
  DFFSRXL imgproc_addr_reg_4_ ( .D(n574), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1306), .QN(n1239) );
  DFFSRXL imgproc_addr_reg_3_ ( .D(n573), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1307), .QN(n1238) );
  DFFSRXL imgproc_addr_reg_2_ ( .D(n572), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1308), .QN(n1237) );
  DFFSRXL imgproc_addr_reg_1_ ( .D(n571), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1309), .QN(n1236) );
  DFFSRXL imgproc_addr_reg_0_ ( .D(n570), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1310), .QN(n1235) );
  DFFSRXL imgproc_addr_reg_7_ ( .D(n577), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1303), .QN(n1242) );
  DFFSRXL col_reg_7_ ( .D(n774), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[7]), 
        .QN(n1259) );
  DFFSRXL imgproc_addr_reg_8_ ( .D(n578), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1302), .QN(n1243) );
  DFFSRXL imgproc_addr_reg_9_ ( .D(n579), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1301), .QN(n1244) );
  DFFSRXL imgproc_addr_reg_10_ ( .D(n580), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1300), .QN(n1245) );
  DFFSRXL imgproc_addr_reg_12_ ( .D(n582), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1298), .QN(n1247) );
  DFFSRXL imgproc_addr_reg_11_ ( .D(n581), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1299), .QN(n1246) );
  DFFSRXL imgproc_addr_reg_13_ ( .D(n583), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1297), .QN(n1248) );
  DFFSRXL imgproc_data_reg_0_ ( .D(n1269), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1318), .QN(n1256) );
  DFFSRXL imgproc_data_reg_1_ ( .D(n1268), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1317), .QN(n1255) );
  DFFSRXL imgproc_data_reg_2_ ( .D(n1267), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1316), .QN(n1254) );
  DFFSRXL imgproc_data_reg_3_ ( .D(n1266), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1315), .QN(n1253) );
  DFFSRXL imgproc_data_reg_4_ ( .D(n1265), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1314), .QN(n1252) );
  DFFSRXL imgproc_data_reg_5_ ( .D(n1264), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1313), .QN(n1251) );
  DFFSRXL imgproc_data_reg_7_ ( .D(n1262), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1311), .QN(n1249) );
  DFFSRXL imgproc_data_reg_6_ ( .D(n1263), .CK(clk), .SN(1'b1), .RN(n12700), 
        .Q(n1312), .QN(n1250) );
  DFFX2 prev_orig_addr_reg_6_ ( .D(n751), .CK(clk), .Q(N672) );
  DFFX2 prev_orig_addr_reg_5_ ( .D(n752), .CK(clk), .Q(N671) );
  DFFX2 prev_orig_addr_reg_4_ ( .D(n753), .CK(clk), .Q(N670) );
  DFFX2 prev_orig_addr_reg_3_ ( .D(n754), .CK(clk), .Q(N669) );
  DFFX2 prev_orig_addr_reg_11_ ( .D(n746), .CK(clk), .Q(n1292) );
  DFFX2 prev_orig_addr_reg_10_ ( .D(n747), .CK(clk), .Q(n1293) );
  DFFX2 prev_orig_addr_reg_8_ ( .D(n749), .CK(clk), .Q(n1295) );
  DFFX2 prev_orig_addr_reg_9_ ( .D(n748), .CK(clk), .Q(n1294) );
  DFFX2 prev_orig_addr_reg_1_ ( .D(n756), .CK(clk), .Q(N165) );
  DFFX2 prev_orig_addr_reg_12_ ( .D(n745), .CK(clk), .Q(n1291), .QN(n912) );
  DFFSRX1 col_reg_0_ ( .D(n781), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[0]), 
        .QN(n1660) );
  DFFX2 prev_orig_addr_reg_13_ ( .D(n744), .CK(clk), .Q(n1290) );
  DFFSRX1 col_reg_2_ ( .D(n779), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[2]), 
        .QN(n1261) );
  DFFSRX1 col_reg_3_ ( .D(n778), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[3]), 
        .QN(n1650) );
  DFFSRX1 col_reg_5_ ( .D(n776), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[5]), 
        .QN(n1257) );
  DFFSRX1 col_reg_1_ ( .D(n780), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[1]), 
        .QN(n1260) );
  DFFSRX1 col_reg_4_ ( .D(n777), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[4]), 
        .QN(n1640) );
  DFFSRX1 col_reg_6_ ( .D(n775), .CK(clk), .SN(1'b1), .RN(n12700), .Q(col[6]), 
        .QN(n1258) );
  DFFX2 array_reg_2__0__0_ ( .D(n655), .CK(clk), .Q(array[106]), .QN(n255) );
  DFFX2 array_reg_0__2__0_ ( .D(n607), .CK(clk), .Q(array[166]), .QN(n1910) );
  DFFX2 array_reg_4__2__0_ ( .D(n735), .CK(clk), .Q(array[14]), .QN(n351) );
  CLKBUFX3 U475 ( .A(N2245), .Y(n792) );
  NAND3X1 U476 ( .A(n1040), .B(n1155), .C(n1214), .Y(n793) );
  AND2X2 U477 ( .A(N1487), .B(add_13_root_add_0_root_add_245_5_carry_17_), .Y(
        n794) );
  AND2X2 U478 ( .A(N1513), .B(N1473), .Y(n797) );
  AND2X2 U479 ( .A(N2126), .B(N1927), .Y(n798) );
  AND2X2 U480 ( .A(N1656), .B(N1351), .Y(n799) );
  AND2X2 U481 ( .A(add_9_root_add_0_root_add_245_5_B_1_), .B(
        add_9_root_add_0_root_add_245_5_A_1_), .Y(n800) );
  AND2X2 U482 ( .A(N2226), .B(N1422), .Y(n801) );
  AND2X2 U483 ( .A(N1634), .B(N1595), .Y(n802) );
  AND2X2 U484 ( .A(N13060), .B(N2072), .Y(n803) );
  AND2X2 U485 ( .A(N1457), .B(N2189), .Y(n804) );
  AND2X2 U486 ( .A(N1620), .B(N2035), .Y(n805) );
  AND2X2 U487 ( .A(N2140), .B(add_7_root_add_0_root_add_245_5_carry_17_), .Y(
        n806) );
  AND2X2 U488 ( .A(N1742), .B(add_6_root_add_0_root_add_245_5_A_3_), .Y(n807)
         );
  AND2X2 U489 ( .A(N1555), .B(N19700), .Y(n808) );
  AND2X2 U490 ( .A(N1389), .B(N1869), .Y(n809) );
  AND2X2 U491 ( .A(N2110), .B(N1321), .Y(n810) );
  AND2X2 U492 ( .A(add_9_root_add_0_root_add_245_5_A_19_), .B(n887), .Y(n811)
         );
  AND2X2 U493 ( .A(N1759), .B(n884), .Y(n812) );
  AND2X2 U494 ( .A(n1291), .B(n908), .Y(n813) );
  NOR4BBX1 U495 ( .AN(n1081), .BN(n1082), .C(n1650), .D(n1640), .Y(n1062) );
  NOR2X1 U496 ( .A(n1260), .B(n1261), .Y(n1081) );
  NOR3XL U497 ( .A(n1660), .B(n1257), .C(n1258), .Y(n1082) );
  AND4XL U498 ( .A(n1257), .B(n1258), .C(n1650), .D(n1640), .Y(n1153) );
  OR3XL U499 ( .A(n1258), .B(n1257), .C(n1650), .Y(n1226) );
  NAND3XL U500 ( .A(n1261), .B(n1153), .C(n1260), .Y(n1074) );
  NAND3XL U501 ( .A(n1153), .B(col[0]), .C(n1260), .Y(n1152) );
  OAI21X2 U502 ( .A0(n942), .A1(n933), .B0(n941), .Y(n1220) );
  OAI21X2 U503 ( .A0(n942), .A1(n1216), .B0(n941), .Y(n1217) );
  OAI21X2 U504 ( .A0(n942), .A1(n1212), .B0(n941), .Y(n1213) );
  OAI21X2 U505 ( .A0(n942), .A1(n932), .B0(n941), .Y(n1211) );
  OAI21X2 U506 ( .A0(n942), .A1(n931), .B0(n941), .Y(n1209) );
  OAI21X2 U507 ( .A0(n942), .A1(n1206), .B0(n941), .Y(n1207) );
  OAI21X2 U508 ( .A0(n942), .A1(n1203), .B0(n941), .Y(n1204) );
  OAI21X2 U509 ( .A0(n942), .A1(n1194), .B0(n941), .Y(n1195) );
  NAND2BXL U510 ( .AN(n1170), .B(n1155), .Y(n1171) );
  OAI21X2 U511 ( .A0(n942), .A1(n943), .B0(n941), .Y(n1222) );
  BUFX4 U512 ( .A(n1170), .Y(n942) );
  INVX12 U513 ( .A(n796), .Y(request) );
  INVX12 U514 ( .A(n795), .Y(imgproc_ready) );
  INVXL U515 ( .A(n848), .Y(n816) );
  INVX12 U516 ( .A(n816), .Y(finish) );
  INVX6 U517 ( .A(rst), .Y(n12700) );
  OAI21X2 U548 ( .A0(n942), .A1(n1197), .B0(n941), .Y(n1198) );
  OAI21X2 U549 ( .A0(n942), .A1(n929), .B0(n941), .Y(n1200) );
  OAI21X2 U550 ( .A0(n942), .A1(n930), .B0(n941), .Y(n1202) );
  OAI21X2 U551 ( .A0(n942), .A1(n1184), .B0(n941), .Y(n1185) );
  BUFX4 U552 ( .A(n1171), .Y(n941) );
  OAI21X2 U553 ( .A0(n942), .A1(n1187), .B0(n941), .Y(n1188) );
  OAI21X2 U554 ( .A0(n942), .A1(n927), .B0(n941), .Y(n1190) );
  OAI21X2 U555 ( .A0(n942), .A1(n928), .B0(n941), .Y(n1192) );
  INVX3 U556 ( .A(n1028), .Y(n1014) );
  NOR2X2 U557 ( .A(n1035), .B(n1039), .Y(n12740) );
  OAI21X2 U558 ( .A0(n942), .A1(n923), .B0(n941), .Y(n1162) );
  AO22X1 U559 ( .A0(n1066), .A1(j[1]), .B0(N179), .B1(n1067), .Y(n772) );
  NOR4BXL U560 ( .AN(j[2]), .B(j[3]), .C(j[1]), .D(j[0]), .Y(n1156) );
  OAI211X4 U561 ( .A0(n1226), .A1(n1227), .B0(n1074), .C0(n1149), .Y(n1027) );
  NOR2X2 U562 ( .A(n1035), .B(n1036), .Y(n12710) );
  OAI21X2 U563 ( .A0(n942), .A1(n924), .B0(n941), .Y(n1175) );
  BUFX12 U564 ( .A(n1312), .Y(imgproc_data[6]) );
  BUFX12 U565 ( .A(n1313), .Y(imgproc_data[5]) );
  BUFX12 U566 ( .A(n1314), .Y(imgproc_data[4]) );
  BUFX12 U567 ( .A(n1315), .Y(imgproc_data[3]) );
  BUFX12 U568 ( .A(n1316), .Y(imgproc_data[2]) );
  BUFX12 U569 ( .A(n1317), .Y(imgproc_data[1]) );
  BUFX12 U570 ( .A(n1318), .Y(imgproc_data[0]) );
  BUFX12 U571 ( .A(n1311), .Y(imgproc_data[7]) );
  NOR2X2 U572 ( .A(n1026), .B(n1062), .Y(n1064) );
  NOR2X2 U573 ( .A(n1043), .B(n1155), .Y(n1223) );
  OAI211X4 U574 ( .A0(n1075), .A1(n1076), .B0(n1049), .C0(n1071), .Y(n1066) );
  NOR2X2 U575 ( .A(n1035), .B(n1037), .Y(n12720) );
  NOR3BX1 U576 ( .AN(n1215), .B(j[0]), .C(j[1]), .Y(n1182) );
  BUFX12 U577 ( .A(n1290), .Y(orig_addr[13]) );
  OAI21X2 U578 ( .A0(n942), .A1(n925), .B0(n941), .Y(n1178) );
  NOR2X2 U579 ( .A(n945), .B(n1048), .Y(n1148) );
  BUFX12 U580 ( .A(n1299), .Y(imgproc_addr[11]) );
  BUFX12 U581 ( .A(n1300), .Y(imgproc_addr[10]) );
  BUFX12 U582 ( .A(n1298), .Y(imgproc_addr[12]) );
  BUFX12 U583 ( .A(n1310), .Y(imgproc_addr[0]) );
  BUFX12 U584 ( .A(n1301), .Y(imgproc_addr[9]) );
  BUFX12 U585 ( .A(n1302), .Y(imgproc_addr[8]) );
  BUFX12 U586 ( .A(n1303), .Y(imgproc_addr[7]) );
  BUFX12 U587 ( .A(n1304), .Y(imgproc_addr[6]) );
  BUFX12 U588 ( .A(n1305), .Y(imgproc_addr[5]) );
  BUFX12 U589 ( .A(n1306), .Y(imgproc_addr[4]) );
  BUFX12 U590 ( .A(n1307), .Y(imgproc_addr[3]) );
  BUFX12 U591 ( .A(n1308), .Y(imgproc_addr[2]) );
  BUFX12 U592 ( .A(n1309), .Y(imgproc_addr[1]) );
  BUFX12 U593 ( .A(n1297), .Y(imgproc_addr[13]) );
  NOR2BX2 U594 ( .AN(n1025), .B(N2238), .Y(n1017) );
  OAI211X4 U595 ( .A0(n1041), .A1(n1076), .B0(n1049), .C0(n1071), .Y(n1077) );
  NOR2X2 U596 ( .A(n1035), .B(n1038), .Y(n12730) );
  NOR3BX1 U597 ( .AN(n1215), .B(n1218), .C(j[1]), .Y(n1179) );
  OA21X2 U598 ( .A0(next_finish), .A1(n1013), .B0(n1048), .Y(n1063) );
  NAND2X2 U599 ( .A(state[0]), .B(n1065), .Y(n1048) );
  BUFX12 U600 ( .A(N165), .Y(orig_addr[1]) );
  OAI21X2 U601 ( .A0(n942), .A1(n926), .B0(n941), .Y(n1181) );
  BUFX12 U602 ( .A(N669), .Y(orig_addr[3]) );
  BUFX12 U603 ( .A(N670), .Y(orig_addr[4]) );
  BUFX12 U604 ( .A(N671), .Y(orig_addr[5]) );
  BUFX12 U605 ( .A(N672), .Y(orig_addr[6]) );
  BUFX12 U606 ( .A(n1294), .Y(orig_addr[9]) );
  BUFX12 U607 ( .A(n1295), .Y(orig_addr[8]) );
  BUFX12 U608 ( .A(n1293), .Y(orig_addr[10]) );
  BUFX12 U609 ( .A(n1292), .Y(orig_addr[11]) );
  INVX12 U610 ( .A(n912), .Y(orig_addr[12]) );
  OAI31X4 U611 ( .A0(n1042), .A1(n1043), .A2(n1044), .B0(n963), .Y(n12750) );
  NOR2BXL U612 ( .AN(n1154), .B(n1041), .Y(n1073) );
  NOR2XL U613 ( .A(n1026), .B(n1027), .Y(n1025) );
  AND2X2 U614 ( .A(n1050), .B(next_imgproc_ready), .Y(n1052) );
  AO22XL U615 ( .A0(n1077), .A1(i[7]), .B0(N163), .B1(n1078), .Y(n758) );
  AO22XL U616 ( .A0(n1066), .A1(j[7]), .B0(N185), .B1(n1067), .Y(n767) );
  AOI22XL U617 ( .A0(N2256), .A1(n1016), .B0(n792), .B1(n1017), .Y(n1018) );
  AND2X2 U618 ( .A(N2238), .B(n1025), .Y(n1016) );
  AND3X2 U619 ( .A(n1071), .B(n1072), .C(n1073), .Y(n1067) );
  AND3X2 U620 ( .A(n1012), .B(n1071), .C(n1041), .Y(n1078) );
  NOR2XL U621 ( .A(n1027), .B(n1151), .Y(n1154) );
  OAI211XL U622 ( .A0(n1047), .A1(n1048), .B0(n1026), .C0(n1049), .Y(n1046) );
  INVXL U623 ( .A(n1027), .Y(n1029) );
  NAND2XL U624 ( .A(n1072), .B(n1027), .Y(n1049) );
  NOR2XL U625 ( .A(n1048), .B(n1027), .Y(n1034) );
  INVXL U626 ( .A(n1048), .Y(n1072) );
  AOI22XL U627 ( .A0(N2254), .A1(n1016), .B0(N2243), .B1(n1017), .Y(n1020) );
  AOI22XL U628 ( .A0(N2255), .A1(n1016), .B0(N2244), .B1(n1017), .Y(n1019) );
  AOI22XL U629 ( .A0(N2252), .A1(n1016), .B0(N2241), .B1(n1017), .Y(n1022) );
  AOI22XL U630 ( .A0(N2253), .A1(n1016), .B0(N2242), .B1(n1017), .Y(n1021) );
  AOI22XL U631 ( .A0(N2250), .A1(n1016), .B0(N2239), .B1(n1017), .Y(n1024) );
  AOI22XL U632 ( .A0(N2251), .A1(n1016), .B0(N2240), .B1(n1017), .Y(n1023) );
  AOI22XL U633 ( .A0(N165), .A1(n921), .B0(N165), .B1(n920), .Y(n1096) );
  AOI22XL U634 ( .A0(N187), .A1(n922), .B0(N165), .B1(n945), .Y(n1095) );
  AOI22XL U635 ( .A0(N192), .A1(n922), .B0(N672), .B1(n945), .Y(n1115) );
  AOI22XL U636 ( .A0(N191), .A1(n922), .B0(N671), .B1(n945), .Y(n1111) );
  AOI22XL U637 ( .A0(N190), .A1(n922), .B0(N670), .B1(n945), .Y(n1107) );
  AOI22XL U638 ( .A0(N189), .A1(n922), .B0(N669), .B1(n945), .Y(n1103) );
  AOI22XL U639 ( .A0(N195), .A1(n922), .B0(orig_addr[9]), .B1(n945), .Y(n1127)
         );
  AOI22XL U640 ( .A0(N194), .A1(n922), .B0(orig_addr[8]), .B1(n945), .Y(n1123)
         );
  AOI22XL U641 ( .A0(N196), .A1(n922), .B0(orig_addr[10]), .B1(n945), .Y(n1131) );
  AOI22XL U642 ( .A0(N197), .A1(n922), .B0(orig_addr[11]), .B1(n945), .Y(n1135) );
  AOI22XL U643 ( .A0(N198), .A1(n922), .B0(n1291), .B1(n945), .Y(n1139) );
  AOI22XL U644 ( .A0(N199), .A1(n922), .B0(n1290), .B1(n945), .Y(n1143) );
  OAI2BB1XL U645 ( .A0N(n1066), .A1N(j[2]), .B0(n1068), .Y(n766) );
  AOI32XL U646 ( .A0(n1069), .A1(n1070), .A2(n1071), .B0(N180), .B1(n1067), 
        .Y(n1068) );
  AO22XL U647 ( .A0(n1077), .A1(i[0]), .B0(N156), .B1(n1078), .Y(n765) );
  AO22XL U648 ( .A0(n1066), .A1(j[0]), .B0(N178), .B1(n1067), .Y(n773) );
  AO22XL U649 ( .A0(n1077), .A1(i[6]), .B0(N162), .B1(n1078), .Y(n759) );
  AO22XL U650 ( .A0(n1077), .A1(i[5]), .B0(N161), .B1(n1078), .Y(n760) );
  AO22XL U651 ( .A0(n1077), .A1(i[4]), .B0(N160), .B1(n1078), .Y(n761) );
  AO22XL U652 ( .A0(n1077), .A1(i[3]), .B0(N159), .B1(n1078), .Y(n762) );
  AO22XL U653 ( .A0(n1077), .A1(i[2]), .B0(N158), .B1(n1078), .Y(n763) );
  AO22XL U654 ( .A0(n1077), .A1(i[1]), .B0(N157), .B1(n1078), .Y(n764) );
  AO22XL U655 ( .A0(n1066), .A1(j[6]), .B0(N184), .B1(n1067), .Y(n768) );
  AO22XL U656 ( .A0(n1066), .A1(j[5]), .B0(N183), .B1(n1067), .Y(n769) );
  AO22XL U657 ( .A0(n1066), .A1(j[4]), .B0(N182), .B1(n1067), .Y(n770) );
  AO22XL U658 ( .A0(n1066), .A1(j[3]), .B0(N181), .B1(n1067), .Y(n771) );
  OR2XL U659 ( .A(N672), .B(sub_203_carry_6_), .Y(sub_203_carry_7_) );
  OR2XL U660 ( .A(N165), .B(n949), .Y(sub_203_carry_2_) );
  OR2XL U661 ( .A(n1292), .B(sub_203_carry_11_), .Y(sub_203_carry_12_) );
  OR2XL U662 ( .A(n1292), .B(sub_139_carry_11_), .Y(sub_139_carry_12_) );
  OR2XL U663 ( .A(n1295), .B(sub_139_carry_8_), .Y(sub_139_carry_9_) );
  OR2XL U664 ( .A(n1294), .B(n892), .Y(sub_203_carry_10_) );
  OR2XL U665 ( .A(n1293), .B(sub_203_carry_10_), .Y(sub_203_carry_11_) );
  OR2XL U666 ( .A(n1293), .B(n893), .Y(sub_139_carry_11_) );
  OR2XL U667 ( .A(N669), .B(sub_203_carry_3_), .Y(sub_203_carry_4_) );
  OR2XL U668 ( .A(N670), .B(sub_203_carry_4_), .Y(sub_203_carry_5_) );
  OR2XL U669 ( .A(N671), .B(sub_203_carry_5_), .Y(sub_203_carry_6_) );
  AND2XL U670 ( .A(N672), .B(n899), .Y(n890) );
  AND2XL U671 ( .A(N165), .B(n949), .Y(n901) );
  AND2XL U672 ( .A(N669), .B(sub_139_carry_3_), .Y(n895) );
  AND2XL U673 ( .A(N670), .B(n895), .Y(n897) );
  AND2XL U674 ( .A(N671), .B(n897), .Y(n899) );
  AND2XL U675 ( .A(n1294), .B(sub_139_carry_9_), .Y(n893) );
  AND2XL U676 ( .A(n1295), .B(sub_203_carry_8_), .Y(n892) );
  OR2XL U677 ( .A(N672), .B(add_146_carry[6]), .Y(add_146_carry[7]) );
  OR2XL U678 ( .A(n1292), .B(r652_carry_11_), .Y(r652_carry_12_) );
  OR2XL U679 ( .A(n1295), .B(r652_carry_8_), .Y(r652_carry_9_) );
  OR2XL U680 ( .A(n1293), .B(n894), .Y(r652_carry_11_) );
  OR2XL U681 ( .A(N669), .B(n947), .Y(add_146_carry[4]) );
  OR2XL U682 ( .A(N670), .B(add_146_carry[4]), .Y(add_146_carry[5]) );
  OR2XL U683 ( .A(N671), .B(add_146_carry[5]), .Y(add_146_carry[6]) );
  AND2XL U684 ( .A(N165), .B(n949), .Y(n902) );
  AND2XL U685 ( .A(N672), .B(n900), .Y(n891) );
  AND2XL U686 ( .A(n1294), .B(n906), .Y(n905) );
  AND2XL U687 ( .A(n1295), .B(n889), .Y(n906) );
  AND2XL U688 ( .A(n1293), .B(n905), .Y(n903) );
  AND2XL U689 ( .A(n1292), .B(n903), .Y(n904) );
  AND2XL U690 ( .A(N669), .B(n888), .Y(n896) );
  AND2XL U691 ( .A(N670), .B(n896), .Y(n898) );
  AND2XL U692 ( .A(N671), .B(n898), .Y(n900) );
  AND2XL U693 ( .A(n1294), .B(r652_carry_9_), .Y(n894) );
  AND2XL U694 ( .A(n1291), .B(n904), .Y(n907) );
  AND2XL U695 ( .A(n1294), .B(n910), .Y(n911) );
  AND2XL U696 ( .A(n1295), .B(n951), .Y(n910) );
  AND2XL U697 ( .A(n1293), .B(n911), .Y(n909) );
  AND2XL U698 ( .A(n1292), .B(n909), .Y(n908) );
  CLKBUFX3 U699 ( .A(n1296), .Y(n951) );
  CLKBUFX3 U700 ( .A(n964), .Y(n961) );
  CLKBUFX3 U701 ( .A(n965), .Y(n959) );
  CLKBUFX3 U702 ( .A(n964), .Y(n960) );
  CLKBUFX3 U703 ( .A(n965), .Y(n958) );
  CLKBUFX3 U704 ( .A(n966), .Y(n956) );
  CLKBUFX3 U705 ( .A(n966), .Y(n957) );
  CLKBUFX3 U706 ( .A(n969), .Y(n963) );
  CLKBUFX3 U707 ( .A(n967), .Y(n962) );
  CLKBUFX3 U708 ( .A(n967), .Y(n954) );
  CLKBUFX3 U709 ( .A(n967), .Y(n955) );
  CLKBUFX3 U710 ( .A(n967), .Y(n953) );
  CLKBUFX3 U711 ( .A(n967), .Y(n952) );
  CLKBUFX3 U712 ( .A(n969), .Y(n964) );
  CLKBUFX3 U713 ( .A(n969), .Y(n965) );
  CLKBUFX3 U714 ( .A(n969), .Y(n966) );
  CLKBUFX3 U715 ( .A(n968), .Y(n967) );
  CLKBUFX3 U716 ( .A(n970), .Y(n969) );
  XOR2X1 U717 ( .A(N2126), .B(N1927), .Y(N1806) );
  XOR2X1 U718 ( .A(N1513), .B(N1473), .Y(
        add_13_root_add_0_root_add_245_5_SUM_3_) );
  XOR2X1 U719 ( .A(N1555), .B(N19700), .Y(add_6_root_add_0_root_add_245_5_A_3_) );
  AND2X2 U720 ( .A(add_9_root_add_0_root_add_245_5_A_15_), .B(
        add_9_root_add_0_root_add_245_5_carry_15_), .Y(n882) );
  AND2X2 U721 ( .A(add_9_root_add_0_root_add_245_5_A_17_), .B(n886), .Y(n883)
         );
  XOR2X1 U722 ( .A(add_9_root_add_0_root_add_245_5_A_15_), .B(
        add_9_root_add_0_root_add_245_5_carry_15_), .Y(N2217) );
  XOR2X1 U723 ( .A(add_9_root_add_0_root_add_245_5_A_17_), .B(n886), .Y(N2219)
         );
  OAI21XL U724 ( .A0(n1214), .A1(n1075), .B0(n1040), .Y(n1170) );
  AND2X2 U725 ( .A(N1758), .B(n885), .Y(n884) );
  XOR2X1 U726 ( .A(N1758), .B(n885), .Y(N1779) );
  AND2X2 U727 ( .A(N1757), .B(add_6_root_add_0_root_add_245_5_carry_18_), .Y(
        n885) );
  XOR2X1 U728 ( .A(N1757), .B(add_6_root_add_0_root_add_245_5_carry_18_), .Y(
        N1778) );
  CLKBUFX3 U729 ( .A(n970), .Y(n968) );
  CLKBUFX3 U730 ( .A(n793), .Y(n970) );
  CLKBUFX3 U731 ( .A(n1093), .Y(n922) );
  AND2XL U732 ( .A(n1148), .B(n1073), .Y(n1093) );
  CLKBUFX3 U733 ( .A(n1090), .Y(n918) );
  AND4XL U734 ( .A(n1148), .B(n1150), .C(n1151), .D(n1029), .Y(n1090) );
  XOR2X1 U735 ( .A(add_9_root_add_0_root_add_245_5_B_1_), .B(
        add_9_root_add_0_root_add_245_5_A_1_), .Y(N2203) );
  XOR2X1 U736 ( .A(N1656), .B(N1351), .Y(N1803) );
  XOR2X1 U737 ( .A(N1595), .B(N1634), .Y(add_9_root_add_0_root_add_245_5_B_1_)
         );
  XOR2X1 U738 ( .A(N1620), .B(N2035), .Y(N1927) );
  XOR2X1 U739 ( .A(N1457), .B(N2189), .Y(N1513) );
  XOR2X1 U740 ( .A(N1742), .B(add_6_root_add_0_root_add_245_5_A_3_), .Y(N1763)
         );
  XOR2X1 U741 ( .A(N2110), .B(N1321), .Y(N19700) );
  XOR2X1 U742 ( .A(N1389), .B(N1869), .Y(N1555) );
  AND2X2 U743 ( .A(add_9_root_add_0_root_add_245_5_A_16_), .B(n882), .Y(n886)
         );
  AND2X2 U744 ( .A(add_9_root_add_0_root_add_245_5_A_18_), .B(n883), .Y(n887)
         );
  XOR2X1 U745 ( .A(N2140), .B(add_7_root_add_0_root_add_245_5_carry_17_), .Y(
        N18200) );
  XOR2X1 U746 ( .A(N1487), .B(add_13_root_add_0_root_add_245_5_carry_17_), .Y(
        add_13_root_add_0_root_add_245_5_SUM_17_) );
  XOR2X1 U747 ( .A(add_9_root_add_0_root_add_245_5_A_16_), .B(n882), .Y(N2218)
         );
  XOR2X1 U748 ( .A(add_9_root_add_0_root_add_245_5_A_18_), .B(n883), .Y(N2220)
         );
  XOR2X1 U749 ( .A(add_9_root_add_0_root_add_245_5_A_19_), .B(n887), .Y(N2221)
         );
  CLKBUFX3 U750 ( .A(n1094), .Y(n945) );
  NAND2X1 U751 ( .A(n1079), .B(n1030), .Y(n1094) );
  XOR2X1 U752 ( .A(N1759), .B(n884), .Y(N17800) );
  CLKBUFX3 U753 ( .A(n1092), .Y(n920) );
  NOR4BBXL U754 ( .AN(n1148), .BN(n1154), .C(n1044), .D(n1155), .Y(n1092) );
  CLKBUFX3 U755 ( .A(n1201), .Y(n930) );
  NAND2XL U756 ( .A(n1182), .B(n1196), .Y(n1201) );
  CLKBUFX3 U757 ( .A(n1199), .Y(n929) );
  NAND2XL U758 ( .A(n1179), .B(n1196), .Y(n1199) );
  CLKBUFX3 U759 ( .A(n1210), .Y(n932) );
  NAND2XL U760 ( .A(n1182), .B(n1205), .Y(n1210) );
  CLKBUFX3 U761 ( .A(n1208), .Y(n931) );
  NAND2XL U762 ( .A(n1179), .B(n1205), .Y(n1208) );
  CLKBUFX3 U763 ( .A(n1219), .Y(n933) );
  NAND2XL U764 ( .A(n1179), .B(n1214), .Y(n1219) );
  CLKINVX1 U765 ( .A(n947), .Y(N166) );
  CLKINVX1 U766 ( .A(n951), .Y(N673) );
  XOR2X1 U767 ( .A(n951), .B(add_146_carry[7]), .Y(N171) );
  CLKBUFX3 U768 ( .A(n1089), .Y(n919) );
  AND4XL U769 ( .A(n1148), .B(n1151), .C(n1029), .D(n1152), .Y(n1089) );
  CLKBUFX3 U770 ( .A(n1091), .Y(n921) );
  AND3XL U771 ( .A(n1154), .B(n1155), .C(n1148), .Y(n1091) );
  CLKBUFX3 U772 ( .A(n1087), .Y(n917) );
  NOR2BXL U773 ( .AN(n1148), .B(n1147), .Y(n1087) );
  CLKBUFX3 U774 ( .A(n1088), .Y(n916) );
  NAND3XL U775 ( .A(n1147), .B(n1027), .C(n1148), .Y(n1088) );
  CLKBUFX3 U776 ( .A(n1221), .Y(n943) );
  NAND2XL U777 ( .A(n1182), .B(n1214), .Y(n1221) );
  CLKBUFX3 U778 ( .A(n1180), .Y(n926) );
  NAND2XL U779 ( .A(n1182), .B(n1173), .Y(n1180) );
  CLKBUFX3 U780 ( .A(n1177), .Y(n925) );
  NAND2XL U781 ( .A(n1179), .B(n1173), .Y(n1177) );
  CLKBUFX3 U782 ( .A(n1191), .Y(n928) );
  NAND2XL U783 ( .A(n1182), .B(n1186), .Y(n1191) );
  CLKBUFX3 U784 ( .A(n1189), .Y(n927) );
  NAND2XL U785 ( .A(n1179), .B(n1186), .Y(n1189) );
  NAND2X2 U786 ( .A(n1176), .B(n1214), .Y(n1216) );
  NAND2X2 U787 ( .A(n1172), .B(n1214), .Y(n1212) );
  NAND2X2 U788 ( .A(n1176), .B(n1186), .Y(n1187) );
  NAND2X2 U789 ( .A(n1172), .B(n1186), .Y(n1184) );
  NAND2X2 U790 ( .A(n1176), .B(n1196), .Y(n1197) );
  NAND2X2 U791 ( .A(n1172), .B(n1196), .Y(n1194) );
  NAND2X2 U792 ( .A(n1176), .B(n1205), .Y(n1206) );
  NAND2X2 U793 ( .A(n1172), .B(n1205), .Y(n1203) );
  CLKBUFX3 U794 ( .A(n1174), .Y(n924) );
  NAND2XL U795 ( .A(n1176), .B(n1173), .Y(n1174) );
  CLKBUFX3 U796 ( .A(n1160), .Y(n923) );
  NAND2XL U797 ( .A(n1172), .B(n1173), .Y(n1160) );
  OR2X1 U798 ( .A(n947), .B(sub_203_carry_2_), .Y(sub_203_carry_3_) );
  OR2X1 U799 ( .A(n951), .B(n890), .Y(sub_139_carry_8_) );
  OR2X1 U800 ( .A(n951), .B(n891), .Y(r652_carry_8_) );
  OR2X1 U801 ( .A(n947), .B(n901), .Y(sub_139_carry_3_) );
  OR2X1 U802 ( .A(n951), .B(sub_203_carry_7_), .Y(sub_203_carry_8_) );
  AND2X2 U803 ( .A(n947), .B(n902), .Y(n888) );
  AND2X2 U804 ( .A(n951), .B(add_146_carry[7]), .Y(n889) );
  XNOR2X1 U805 ( .A(n951), .B(sub_203_carry_7_), .Y(N1002) );
  XNOR2X1 U806 ( .A(n951), .B(n891), .Y(N134) );
  XNOR2X1 U807 ( .A(n951), .B(n890), .Y(N120) );
  CLKAND2X3 U808 ( .A(n1031), .B(n1048), .Y(n1233) );
  AND2X2 U809 ( .A(n1233), .B(n1069), .Y(n1234) );
  XNOR2X1 U810 ( .A(n947), .B(sub_203_carry_2_), .Y(N997) );
  XNOR2X1 U811 ( .A(n947), .B(n901), .Y(N115) );
  XOR2X1 U812 ( .A(n947), .B(n902), .Y(N129) );
  AND2X2 U813 ( .A(n1060), .B(n1048), .Y(n1050) );
  XOR2X1 U814 ( .A(N13060), .B(N2072), .Y(N1634) );
  XOR2X1 U815 ( .A(N2226), .B(N1422), .Y(N1595) );
  CLKBUFX3 U816 ( .A(n1161), .Y(n934) );
  NAND2XL U817 ( .A(orig_data[0]), .B(n1223), .Y(n1161) );
  CLKBUFX3 U818 ( .A(n1163), .Y(n935) );
  NAND2XL U819 ( .A(orig_data[1]), .B(n1223), .Y(n1163) );
  CLKBUFX3 U820 ( .A(n1164), .Y(n936) );
  NAND2XL U821 ( .A(orig_data[2]), .B(n1223), .Y(n1164) );
  CLKBUFX3 U822 ( .A(n1165), .Y(n937) );
  NAND2XL U823 ( .A(orig_data[3]), .B(n1223), .Y(n1165) );
  CLKBUFX3 U824 ( .A(n1166), .Y(n938) );
  NAND2XL U825 ( .A(orig_data[4]), .B(n1223), .Y(n1166) );
  CLKBUFX3 U826 ( .A(n1167), .Y(n939) );
  NAND2XL U827 ( .A(orig_data[5]), .B(n1223), .Y(n1167) );
  CLKBUFX3 U828 ( .A(n1168), .Y(n940) );
  NAND2XL U829 ( .A(orig_data[6]), .B(n1223), .Y(n1168) );
  CLKBUFX3 U830 ( .A(n1169), .Y(n944) );
  NAND2XL U831 ( .A(orig_data[7]), .B(n1223), .Y(n1169) );
  XNOR2XL U832 ( .A(N672), .B(add_146_carry[6]), .Y(N170) );
  XNOR2XL U833 ( .A(N671), .B(add_146_carry[5]), .Y(N169) );
  XNOR2XL U834 ( .A(N670), .B(add_146_carry[4]), .Y(N168) );
  XNOR2XL U835 ( .A(N669), .B(n947), .Y(N167) );
  XOR2XL U836 ( .A(n1295), .B(n951), .Y(N674) );
  XOR2XL U837 ( .A(n1295), .B(n889), .Y(N172) );
  XOR2XL U838 ( .A(n1294), .B(n910), .Y(N675) );
  XOR2XL U839 ( .A(n1294), .B(n906), .Y(N173) );
  XOR2XL U840 ( .A(n1293), .B(n911), .Y(N676) );
  XOR2XL U841 ( .A(n1293), .B(n905), .Y(N174) );
  XOR2XL U842 ( .A(n1292), .B(n909), .Y(N677) );
  XOR2XL U843 ( .A(n1292), .B(n903), .Y(N175) );
  XOR2XL U844 ( .A(n1291), .B(n908), .Y(N678) );
  XOR2XL U845 ( .A(n1291), .B(n904), .Y(N176) );
  XOR2XL U846 ( .A(n1290), .B(n813), .Y(N679) );
  XOR2XL U847 ( .A(n1290), .B(n907), .Y(N177) );
  XNOR2XL U848 ( .A(n1291), .B(sub_139_carry_12_), .Y(N125) );
  XNOR2XL U849 ( .A(n1290), .B(r652_carry_13_), .Y(N140) );
  NAND2X1 U850 ( .A(n912), .B(n915), .Y(r652_carry_13_) );
  CLKINVX1 U851 ( .A(r652_carry_12_), .Y(n915) );
  XNOR2XL U852 ( .A(n1290), .B(sub_203_carry_13_), .Y(N1008) );
  NAND2X1 U853 ( .A(n912), .B(n913), .Y(sub_203_carry_13_) );
  CLKINVX1 U854 ( .A(sub_203_carry_12_), .Y(n913) );
  XNOR2XL U855 ( .A(n1290), .B(sub_139_carry_13_), .Y(N126) );
  NAND2X1 U856 ( .A(n912), .B(n914), .Y(sub_139_carry_13_) );
  CLKINVX1 U857 ( .A(sub_139_carry_12_), .Y(n914) );
  XNOR2XL U858 ( .A(n1293), .B(n894), .Y(N137) );
  XNOR2XL U859 ( .A(n1292), .B(r652_carry_11_), .Y(N138) );
  XNOR2XL U860 ( .A(n1291), .B(r652_carry_12_), .Y(N139) );
  XNOR2XL U861 ( .A(n1295), .B(r652_carry_8_), .Y(N135) );
  XNOR2XL U862 ( .A(n1293), .B(n893), .Y(N123) );
  XNOR2XL U863 ( .A(n1292), .B(sub_139_carry_11_), .Y(N124) );
  XNOR2XL U864 ( .A(n1295), .B(sub_139_carry_8_), .Y(N121) );
  XNOR2XL U865 ( .A(n1293), .B(sub_203_carry_10_), .Y(N1005) );
  XNOR2XL U866 ( .A(n1292), .B(sub_203_carry_11_), .Y(N1006) );
  XNOR2XL U867 ( .A(n1291), .B(sub_203_carry_12_), .Y(N1007) );
  XNOR2XL U868 ( .A(n1294), .B(n892), .Y(N1004) );
  XOR2XL U869 ( .A(n1294), .B(r652_carry_9_), .Y(N136) );
  XOR2XL U870 ( .A(n1294), .B(sub_139_carry_9_), .Y(N122) );
  XOR2XL U871 ( .A(n1295), .B(sub_203_carry_8_), .Y(N1003) );
  XNOR2XL U872 ( .A(N672), .B(sub_203_carry_6_), .Y(N1001) );
  XNOR2XL U873 ( .A(N671), .B(sub_203_carry_5_), .Y(N1000) );
  XNOR2XL U874 ( .A(N670), .B(sub_203_carry_4_), .Y(N999) );
  XOR2XL U875 ( .A(N672), .B(n900), .Y(N133) );
  XOR2XL U876 ( .A(N671), .B(n898), .Y(N132) );
  XOR2XL U877 ( .A(N670), .B(n896), .Y(N131) );
  XOR2XL U878 ( .A(N672), .B(n899), .Y(N119) );
  XOR2XL U879 ( .A(N671), .B(n897), .Y(N118) );
  XOR2XL U880 ( .A(N670), .B(n895), .Y(N117) );
  CLKBUFX3 U881 ( .A(N668), .Y(n947) );
  CLKBUFX3 U882 ( .A(N164), .Y(n949) );
  XNOR2XL U883 ( .A(N669), .B(sub_203_carry_3_), .Y(N998) );
  XNOR2XL U884 ( .A(N165), .B(n949), .Y(N996) );
  XOR2XL U885 ( .A(N669), .B(n888), .Y(N130) );
  XOR2XL U886 ( .A(N669), .B(sub_139_carry_3_), .Y(N116) );
  XOR2XL U887 ( .A(N165), .B(n949), .Y(N128) );
  XOR2XL U888 ( .A(N165), .B(n949), .Y(N114) );
  BUFX12 U889 ( .A(N164), .Y(orig_addr[0]) );
  BUFX12 U890 ( .A(N668), .Y(orig_addr[2]) );
  BUFX12 U891 ( .A(n1296), .Y(orig_addr[7]) );
  CLKBUFX3 U892 ( .A(n12700), .Y(n971) );
  XNOR2X1 U893 ( .A(array[141]), .B(mult_242_2_n3), .Y(N1507) );
  NOR2X1 U894 ( .A(mult_242_2_n3), .B(array[141]), .Y(n972) );
  XNOR2X1 U895 ( .A(n980), .B(n972), .Y(N1508) );
  NAND2X1 U896 ( .A(n972), .B(n980), .Y(n973) );
  XNOR2X1 U897 ( .A(array[143]), .B(n973), .Y(N1509) );
  XNOR2X1 U898 ( .A(array[126]), .B(mult_242_4_n3), .Y(N1591) );
  NOR2X1 U899 ( .A(mult_242_4_n3), .B(array[126]), .Y(n982) );
  XNOR2X1 U900 ( .A(n990), .B(n982), .Y(N1592) );
  NAND2X1 U901 ( .A(n982), .B(n990), .Y(n983) );
  XNOR2X1 U902 ( .A(array[128]), .B(n983), .Y(N1593) );
  XNOR2X1 U903 ( .A(array[63]), .B(mult_244_2_n3), .Y(N1921) );
  NOR2X1 U904 ( .A(mult_244_2_n3), .B(array[63]), .Y(n992) );
  XNOR2X1 U905 ( .A(n10000), .B(n992), .Y(N1922) );
  NAND2X1 U906 ( .A(n992), .B(n10000), .Y(n993) );
  XNOR2X1 U907 ( .A(array[65]), .B(n993), .Y(N1923) );
  XNOR2X1 U908 ( .A(array[48]), .B(mult_244_4_n3), .Y(N2006) );
  NOR2X1 U909 ( .A(mult_244_4_n3), .B(array[48]), .Y(n10020) );
  XNOR2X1 U910 ( .A(n1010), .B(n10020), .Y(N2007) );
  NAND2X1 U911 ( .A(n10020), .B(n1010), .Y(n10030) );
  XNOR2X1 U912 ( .A(array[50]), .B(n10030), .Y(N2008) );
  CLKINVX1 U913 ( .A(n949), .Y(N127) );
  OAI2BB1X1 U914 ( .A0N(n1012), .A1N(orig_ready), .B0(n1013), .Y(next_request)
         );
  OAI21XL U915 ( .A0(n1249), .A1(n1014), .B0(n1015), .Y(n1262) );
  AOI22X1 U916 ( .A0(N2257), .A1(n1016), .B0(N2246), .B1(n1017), .Y(n1015) );
  OAI21XL U917 ( .A0(n1250), .A1(n1014), .B0(n1018), .Y(n1263) );
  OAI21XL U918 ( .A0(n1251), .A1(n1014), .B0(n1019), .Y(n1264) );
  OAI21XL U919 ( .A0(n1252), .A1(n1014), .B0(n1020), .Y(n1265) );
  OAI21XL U920 ( .A0(n1253), .A1(n1014), .B0(n1021), .Y(n1266) );
  OAI21XL U921 ( .A0(n1254), .A1(n1014), .B0(n1022), .Y(n1267) );
  OAI21XL U922 ( .A0(n1255), .A1(n1014), .B0(n1023), .Y(n1268) );
  OAI21XL U923 ( .A0(n1256), .A1(n1014), .B0(n1024), .Y(n1269) );
  OAI211X1 U924 ( .A0(n1029), .A1(n1030), .B0(n1031), .C0(n1032), .Y(n1028) );
  NOR2X1 U925 ( .A(n1033), .B(n1034), .Y(n1032) );
  NAND2X1 U926 ( .A(n1040), .B(n1041), .Y(n1035) );
  NAND4BX1 U927 ( .AN(n1033), .B(n1013), .C(n1045), .D(n1026), .Y(n791) );
  NOR2BX1 U928 ( .AN(n1046), .B(n1033), .Y(n790) );
  OAI2BB2XL U929 ( .B0(n1050), .B1(n1051), .A0N(N1270), .A1N(n1052), .Y(n789)
         );
  OAI2BB2XL U930 ( .B0(n1050), .B1(n1053), .A0N(N1271), .A1N(n1052), .Y(n788)
         );
  OAI2BB2XL U931 ( .B0(n1050), .B1(n1054), .A0N(N1272), .A1N(n1052), .Y(n787)
         );
  OAI2BB2XL U932 ( .B0(n1050), .B1(n1055), .A0N(N1273), .A1N(n1052), .Y(n786)
         );
  OAI2BB2XL U933 ( .B0(n1050), .B1(n1056), .A0N(N1274), .A1N(n1052), .Y(n785)
         );
  OAI2BB2XL U934 ( .B0(n1050), .B1(n1057), .A0N(N1275), .A1N(n1052), .Y(n784)
         );
  OAI2BB2XL U935 ( .B0(n1050), .B1(n1058), .A0N(N1276), .A1N(n1052), .Y(n783)
         );
  OAI2BB2XL U936 ( .B0(n1050), .B1(n1059), .A0N(N1277), .A1N(n1052), .Y(n782)
         );
  OAI2BB2XL U937 ( .B0(n1061), .B1(n1059), .A0N(n1013), .A1N(n1062), .Y(n1060)
         );
  OAI2BB2XL U938 ( .B0(n1660), .B1(n1063), .A0N(N1282), .A1N(n1064), .Y(n781)
         );
  OAI2BB2XL U939 ( .B0(n1260), .B1(n1063), .A0N(N1283), .A1N(n1064), .Y(n780)
         );
  OAI2BB2XL U940 ( .B0(n1261), .B1(n1063), .A0N(N1284), .A1N(n1064), .Y(n779)
         );
  OAI2BB2XL U941 ( .B0(n1650), .B1(n1063), .A0N(N1285), .A1N(n1064), .Y(n778)
         );
  OAI2BB2XL U942 ( .B0(n1640), .B1(n1063), .A0N(N1286), .A1N(n1064), .Y(n777)
         );
  OAI2BB2XL U943 ( .B0(n1257), .B1(n1063), .A0N(N1287), .A1N(n1064), .Y(n776)
         );
  OAI2BB2XL U944 ( .B0(n1258), .B1(n1063), .A0N(N1288), .A1N(n1064), .Y(n775)
         );
  OAI2BB2XL U945 ( .B0(n1259), .B1(n1063), .A0N(N1289), .A1N(n1064), .Y(n774)
         );
  CLKINVX1 U946 ( .A(next_imgproc_ready), .Y(n1026) );
  NOR2X1 U947 ( .A(n1030), .B(row[7]), .Y(next_imgproc_ready) );
  AOI21X1 U948 ( .A0(state[0]), .A1(state[1]), .B0(n1061), .Y(n1013) );
  NOR2X1 U949 ( .A(n1059), .B(n1065), .Y(next_finish) );
  OAI21XL U950 ( .A0(n1074), .A1(col[0]), .B0(n1075), .Y(n1070) );
  CLKINVX1 U951 ( .A(n1045), .Y(n1012) );
  NAND2X1 U952 ( .A(n1034), .B(n1047), .Y(n1045) );
  AND2X1 U953 ( .A(n1079), .B(n1080), .Y(n1071) );
  OAI21XL U954 ( .A0(n1062), .A1(row[7]), .B0(n1069), .Y(n1080) );
  NAND2X1 U955 ( .A(n1072), .B(n1047), .Y(n1076) );
  NAND4X1 U956 ( .A(n1083), .B(n1084), .C(n1085), .D(n1086), .Y(n757) );
  AOI2BB2X1 U957 ( .B0(N127), .B1(n917), .A0N(n1660), .A1N(n916), .Y(n1086) );
  AOI22X1 U958 ( .A0(N127), .A1(n919), .B0(N127), .B1(n918), .Y(n1085) );
  AOI22X1 U959 ( .A0(n949), .A1(n921), .B0(n949), .B1(n920), .Y(n1084) );
  AOI22X1 U960 ( .A0(N186), .A1(n922), .B0(n949), .B1(n945), .Y(n1083) );
  NAND4X1 U961 ( .A(n1095), .B(n1096), .C(n1097), .D(n1098), .Y(n756) );
  AOI2BB2X1 U962 ( .B0(N996), .B1(n917), .A0N(n1260), .A1N(n916), .Y(n1098) );
  AOI22X1 U963 ( .A0(N128), .A1(n919), .B0(N114), .B1(n918), .Y(n1097) );
  NAND4X1 U964 ( .A(n1099), .B(n1100), .C(n1101), .D(n1102), .Y(n755) );
  AOI2BB2X1 U965 ( .B0(N997), .B1(n917), .A0N(n1261), .A1N(n916), .Y(n1102) );
  AOI22X1 U966 ( .A0(N129), .A1(n919), .B0(N115), .B1(n918), .Y(n1101) );
  AOI22X1 U967 ( .A0(n947), .A1(n921), .B0(N166), .B1(n920), .Y(n1100) );
  AOI22X1 U968 ( .A0(N188), .A1(n922), .B0(n947), .B1(n945), .Y(n1099) );
  NAND4X1 U969 ( .A(n1103), .B(n1104), .C(n1105), .D(n1106), .Y(n754) );
  AOI2BB2X1 U970 ( .B0(N998), .B1(n917), .A0N(n1650), .A1N(n916), .Y(n1106) );
  AOI22X1 U971 ( .A0(N130), .A1(n919), .B0(N116), .B1(n918), .Y(n1105) );
  AOI22X1 U972 ( .A0(N669), .A1(n921), .B0(N167), .B1(n920), .Y(n1104) );
  NAND4X1 U973 ( .A(n1107), .B(n1108), .C(n1109), .D(n1110), .Y(n753) );
  AOI2BB2X1 U974 ( .B0(N999), .B1(n917), .A0N(n1640), .A1N(n916), .Y(n1110) );
  AOI22X1 U975 ( .A0(N131), .A1(n919), .B0(N117), .B1(n918), .Y(n1109) );
  AOI22X1 U976 ( .A0(N670), .A1(n921), .B0(N168), .B1(n920), .Y(n1108) );
  NAND4X1 U977 ( .A(n1111), .B(n1112), .C(n1113), .D(n1114), .Y(n752) );
  AOI2BB2X1 U978 ( .B0(N1000), .B1(n917), .A0N(n1257), .A1N(n916), .Y(n1114)
         );
  AOI22X1 U979 ( .A0(N132), .A1(n919), .B0(N118), .B1(n918), .Y(n1113) );
  AOI22X1 U980 ( .A0(N671), .A1(n921), .B0(N169), .B1(n920), .Y(n1112) );
  NAND4X1 U981 ( .A(n1115), .B(n1116), .C(n1117), .D(n1118), .Y(n751) );
  AOI2BB2X1 U982 ( .B0(N1001), .B1(n917), .A0N(n1258), .A1N(n916), .Y(n1118)
         );
  AOI22X1 U983 ( .A0(N133), .A1(n919), .B0(N119), .B1(n918), .Y(n1117) );
  AOI22X1 U984 ( .A0(N672), .A1(n921), .B0(N170), .B1(n920), .Y(n1116) );
  NAND4X1 U985 ( .A(n1119), .B(n1120), .C(n1121), .D(n1122), .Y(n750) );
  AOI2BB2X1 U986 ( .B0(N1002), .B1(n917), .A0N(n1051), .A1N(n916), .Y(n1122)
         );
  AOI22X1 U987 ( .A0(N134), .A1(n919), .B0(N120), .B1(n918), .Y(n1121) );
  AOI22X1 U988 ( .A0(N673), .A1(n921), .B0(N171), .B1(n920), .Y(n1120) );
  AOI22X1 U989 ( .A0(N193), .A1(n922), .B0(n951), .B1(n945), .Y(n1119) );
  NAND4X1 U990 ( .A(n1123), .B(n1124), .C(n1125), .D(n1126), .Y(n749) );
  AOI2BB2X1 U991 ( .B0(N1003), .B1(n917), .A0N(n1053), .A1N(n916), .Y(n1126)
         );
  AOI22X1 U992 ( .A0(N135), .A1(n919), .B0(N121), .B1(n918), .Y(n1125) );
  AOI22X1 U993 ( .A0(N674), .A1(n921), .B0(N172), .B1(n920), .Y(n1124) );
  NAND4X1 U994 ( .A(n1127), .B(n1128), .C(n1129), .D(n1130), .Y(n748) );
  AOI2BB2X1 U995 ( .B0(N1004), .B1(n917), .A0N(n1054), .A1N(n916), .Y(n1130)
         );
  AOI22X1 U996 ( .A0(N136), .A1(n919), .B0(N122), .B1(n918), .Y(n1129) );
  AOI22X1 U997 ( .A0(N675), .A1(n921), .B0(N173), .B1(n920), .Y(n1128) );
  NAND4X1 U998 ( .A(n1131), .B(n1132), .C(n1133), .D(n1134), .Y(n747) );
  AOI2BB2X1 U999 ( .B0(N1005), .B1(n917), .A0N(n1055), .A1N(n916), .Y(n1134)
         );
  AOI22X1 U1000 ( .A0(N137), .A1(n919), .B0(N123), .B1(n918), .Y(n1133) );
  AOI22X1 U1001 ( .A0(N676), .A1(n921), .B0(N174), .B1(n920), .Y(n1132) );
  NAND4X1 U1002 ( .A(n1135), .B(n1136), .C(n1137), .D(n1138), .Y(n746) );
  AOI2BB2X1 U1003 ( .B0(N1006), .B1(n917), .A0N(n1056), .A1N(n916), .Y(n1138)
         );
  AOI22X1 U1004 ( .A0(N138), .A1(n919), .B0(N124), .B1(n918), .Y(n1137) );
  AOI22X1 U1005 ( .A0(N677), .A1(n921), .B0(N175), .B1(n920), .Y(n1136) );
  NAND4X1 U1006 ( .A(n1139), .B(n1140), .C(n1141), .D(n1142), .Y(n745) );
  AOI2BB2X1 U1007 ( .B0(N1007), .B1(n917), .A0N(n1057), .A1N(n916), .Y(n1142)
         );
  AOI22X1 U1008 ( .A0(N139), .A1(n919), .B0(N125), .B1(n918), .Y(n1141) );
  AOI22X1 U1009 ( .A0(N678), .A1(n921), .B0(N176), .B1(n920), .Y(n1140) );
  NAND4X1 U1010 ( .A(n1143), .B(n1144), .C(n1145), .D(n1146), .Y(n744) );
  AOI2BB2X1 U1011 ( .B0(N1008), .B1(n917), .A0N(n1058), .A1N(n916), .Y(n1146)
         );
  NAND3X1 U1012 ( .A(n1149), .B(n1261), .C(n1150), .Y(n1147) );
  AOI22X1 U1013 ( .A0(N140), .A1(n919), .B0(N126), .B1(n918), .Y(n1145) );
  CLKINVX1 U1014 ( .A(n1152), .Y(n1150) );
  AOI22X1 U1015 ( .A0(N679), .A1(n921), .B0(N177), .B1(n920), .Y(n1144) );
  NAND2X1 U1016 ( .A(n1075), .B(n1044), .Y(n1041) );
  NAND2X1 U1017 ( .A(n1156), .B(n1157), .Y(n1044) );
  NOR4X1 U1018 ( .A(j[7]), .B(j[6]), .C(j[5]), .D(j[4]), .Y(n1157) );
  CLKINVX1 U1019 ( .A(n1047), .Y(n1151) );
  NAND4X1 U1020 ( .A(i[2]), .B(i[0]), .C(n1158), .D(n1159), .Y(n1047) );
  OAI222XL U1021 ( .A0(n923), .A1(n934), .B0(n359), .B1(n1162), .C0(n367), 
        .C1(n963), .Y(n743) );
  OAI222XL U1022 ( .A0(n923), .A1(n935), .B0(n358), .B1(n1162), .C0(n366), 
        .C1(n963), .Y(n742) );
  OAI222XL U1023 ( .A0(n923), .A1(n936), .B0(n357), .B1(n1162), .C0(n365), 
        .C1(n963), .Y(n741) );
  OAI222XL U1024 ( .A0(n923), .A1(n937), .B0(n356), .B1(n1162), .C0(n364), 
        .C1(n963), .Y(n740) );
  OAI222XL U1025 ( .A0(n923), .A1(n938), .B0(n355), .B1(n1162), .C0(n363), 
        .C1(n962), .Y(n739) );
  OAI222XL U1026 ( .A0(n923), .A1(n939), .B0(n354), .B1(n1162), .C0(n362), 
        .C1(n962), .Y(n738) );
  OAI222XL U1027 ( .A0(n923), .A1(n940), .B0(n353), .B1(n1162), .C0(n361), 
        .C1(n962), .Y(n737) );
  OAI222XL U1028 ( .A0(n923), .A1(n944), .B0(n352), .B1(n1162), .C0(n360), 
        .C1(n962), .Y(n736) );
  OAI222XL U1029 ( .A0(n934), .A1(n924), .B0(n351), .B1(n1175), .C0(n359), 
        .C1(n962), .Y(n735) );
  OAI222XL U1030 ( .A0(n935), .A1(n924), .B0(n350), .B1(n1175), .C0(n358), 
        .C1(n962), .Y(n734) );
  OAI222XL U1031 ( .A0(n936), .A1(n924), .B0(n349), .B1(n1175), .C0(n357), 
        .C1(n962), .Y(n733) );
  OAI222XL U1032 ( .A0(n937), .A1(n924), .B0(n348), .B1(n1175), .C0(n356), 
        .C1(n962), .Y(n732) );
  OAI222XL U1033 ( .A0(n938), .A1(n924), .B0(n347), .B1(n1175), .C0(n355), 
        .C1(n962), .Y(n731) );
  OAI222XL U1034 ( .A0(n939), .A1(n924), .B0(n346), .B1(n1175), .C0(n354), 
        .C1(n962), .Y(n730) );
  OAI222XL U1035 ( .A0(n940), .A1(n924), .B0(n345), .B1(n1175), .C0(n353), 
        .C1(n962), .Y(n729) );
  OAI222XL U1036 ( .A0(n944), .A1(n924), .B0(n344), .B1(n1175), .C0(n352), 
        .C1(n962), .Y(n728) );
  OAI222XL U1037 ( .A0(n934), .A1(n925), .B0(n343), .B1(n1178), .C0(n351), 
        .C1(n962), .Y(n727) );
  OAI222XL U1038 ( .A0(n935), .A1(n925), .B0(n342), .B1(n1178), .C0(n350), 
        .C1(n961), .Y(n726) );
  OAI222XL U1039 ( .A0(n936), .A1(n925), .B0(n341), .B1(n1178), .C0(n349), 
        .C1(n961), .Y(n725) );
  OAI222XL U1040 ( .A0(n937), .A1(n925), .B0(n340), .B1(n1178), .C0(n348), 
        .C1(n961), .Y(n724) );
  OAI222XL U1041 ( .A0(n938), .A1(n925), .B0(n339), .B1(n1178), .C0(n347), 
        .C1(n961), .Y(n723) );
  OAI222XL U1042 ( .A0(n939), .A1(n925), .B0(n338), .B1(n1178), .C0(n346), 
        .C1(n961), .Y(n722) );
  OAI222XL U1043 ( .A0(n940), .A1(n925), .B0(n337), .B1(n1178), .C0(n345), 
        .C1(n961), .Y(n721) );
  OAI222XL U1044 ( .A0(n944), .A1(n925), .B0(n336), .B1(n1178), .C0(n344), 
        .C1(n961), .Y(n720) );
  OAI222XL U1045 ( .A0(n934), .A1(n926), .B0(n335), .B1(n1181), .C0(n343), 
        .C1(n961), .Y(n719) );
  OAI222XL U1046 ( .A0(n935), .A1(n926), .B0(n334), .B1(n1181), .C0(n342), 
        .C1(n961), .Y(n718) );
  OAI222XL U1047 ( .A0(n936), .A1(n926), .B0(n333), .B1(n1181), .C0(n341), 
        .C1(n961), .Y(n717) );
  OAI222XL U1048 ( .A0(n937), .A1(n926), .B0(n332), .B1(n1181), .C0(n340), 
        .C1(n961), .Y(n716) );
  OAI222XL U1049 ( .A0(n938), .A1(n926), .B0(n331), .B1(n1181), .C0(n339), 
        .C1(n961), .Y(n715) );
  OAI222XL U1050 ( .A0(n939), .A1(n926), .B0(n330), .B1(n1181), .C0(n338), 
        .C1(n961), .Y(n714) );
  OAI222XL U1051 ( .A0(n940), .A1(n926), .B0(n329), .B1(n1181), .C0(n337), 
        .C1(n960), .Y(n713) );
  OAI222XL U1052 ( .A0(n944), .A1(n926), .B0(n328), .B1(n1181), .C0(n336), 
        .C1(n960), .Y(n712) );
  CLKINVX1 U1053 ( .A(n1036), .Y(n1173) );
  NAND4X1 U1054 ( .A(i[2]), .B(n1158), .C(n1183), .D(n1159), .Y(n1036) );
  OAI222XL U1055 ( .A0(n934), .A1(n1184), .B0(n10040), .B1(n1185), .C0(n327), 
        .C1(n960), .Y(n711) );
  OAI222XL U1056 ( .A0(n935), .A1(n1184), .B0(n10050), .B1(n1185), .C0(n326), 
        .C1(n960), .Y(n710) );
  OAI222XL U1057 ( .A0(n936), .A1(n1184), .B0(n10060), .B1(n1185), .C0(n325), 
        .C1(n960), .Y(n709) );
  OAI222XL U1058 ( .A0(n937), .A1(n1184), .B0(n10070), .B1(n1185), .C0(n324), 
        .C1(n960), .Y(n708) );
  OAI222XL U1059 ( .A0(n938), .A1(n1184), .B0(n10080), .B1(n1185), .C0(n323), 
        .C1(n960), .Y(n707) );
  OAI222XL U1060 ( .A0(n939), .A1(n1184), .B0(n1009), .B1(n1185), .C0(n322), 
        .C1(n960), .Y(n706) );
  OAI222XL U1061 ( .A0(n940), .A1(n1184), .B0(n1010), .B1(n1185), .C0(n321), 
        .C1(n960), .Y(n705) );
  OAI222XL U1062 ( .A0(n944), .A1(n1184), .B0(n1011), .B1(n1185), .C0(n320), 
        .C1(n960), .Y(n704) );
  OAI222XL U1063 ( .A0(n934), .A1(n1187), .B0(n311), .B1(n1188), .C0(n10040), 
        .C1(n960), .Y(n703) );
  OAI222XL U1064 ( .A0(n935), .A1(n1187), .B0(n310), .B1(n1188), .C0(n10050), 
        .C1(n960), .Y(n702) );
  OAI222XL U1065 ( .A0(n936), .A1(n1187), .B0(n309), .B1(n1188), .C0(n10060), 
        .C1(n960), .Y(n701) );
  OAI222XL U1066 ( .A0(n937), .A1(n1187), .B0(n308), .B1(n1188), .C0(n10070), 
        .C1(n959), .Y(n700) );
  OAI222XL U1067 ( .A0(n938), .A1(n1187), .B0(n307), .B1(n1188), .C0(n10080), 
        .C1(n959), .Y(n699) );
  OAI222XL U1068 ( .A0(n939), .A1(n1187), .B0(n306), .B1(n1188), .C0(n1009), 
        .C1(n959), .Y(n698) );
  OAI222XL U1069 ( .A0(n940), .A1(n1187), .B0(n305), .B1(n1188), .C0(n1010), 
        .C1(n959), .Y(n697) );
  OAI222XL U1070 ( .A0(n944), .A1(n1187), .B0(n304), .B1(n1188), .C0(n1011), 
        .C1(n959), .Y(n696) );
  OAI222XL U1071 ( .A0(n934), .A1(n927), .B0(n994), .B1(n1190), .C0(n311), 
        .C1(n959), .Y(n695) );
  OAI222XL U1072 ( .A0(n935), .A1(n927), .B0(n995), .B1(n1190), .C0(n310), 
        .C1(n959), .Y(n694) );
  OAI222XL U1073 ( .A0(n936), .A1(n927), .B0(n9960), .B1(n1190), .C0(n309), 
        .C1(n959), .Y(n693) );
  OAI222XL U1074 ( .A0(n937), .A1(n927), .B0(n9970), .B1(n1190), .C0(n308), 
        .C1(n959), .Y(n692) );
  OAI222XL U1075 ( .A0(n938), .A1(n927), .B0(n9980), .B1(n1190), .C0(n307), 
        .C1(n959), .Y(n691) );
  OAI222XL U1076 ( .A0(n939), .A1(n927), .B0(n9990), .B1(n1190), .C0(n306), 
        .C1(n959), .Y(n690) );
  OAI222XL U1077 ( .A0(n940), .A1(n927), .B0(n10000), .B1(n1190), .C0(n305), 
        .C1(n959), .Y(n689) );
  OAI222XL U1078 ( .A0(n944), .A1(n927), .B0(n10010), .B1(n1190), .C0(n304), 
        .C1(n959), .Y(n688) );
  OAI222XL U1079 ( .A0(n934), .A1(n928), .B0(n295), .B1(n1192), .C0(n994), 
        .C1(n958), .Y(n687) );
  OAI222XL U1080 ( .A0(n935), .A1(n928), .B0(n294), .B1(n1192), .C0(n995), 
        .C1(n958), .Y(n686) );
  OAI222XL U1081 ( .A0(n936), .A1(n928), .B0(n293), .B1(n1192), .C0(n9960), 
        .C1(n958), .Y(n685) );
  OAI222XL U1082 ( .A0(n937), .A1(n928), .B0(n292), .B1(n1192), .C0(n9970), 
        .C1(n958), .Y(n684) );
  OAI222XL U1083 ( .A0(n938), .A1(n928), .B0(n291), .B1(n1192), .C0(n9980), 
        .C1(n958), .Y(n683) );
  OAI222XL U1084 ( .A0(n939), .A1(n928), .B0(n290), .B1(n1192), .C0(n9990), 
        .C1(n958), .Y(n682) );
  OAI222XL U1085 ( .A0(n940), .A1(n928), .B0(n289), .B1(n1192), .C0(n10000), 
        .C1(n958), .Y(n681) );
  OAI222XL U1086 ( .A0(n944), .A1(n928), .B0(n288), .B1(n1192), .C0(n10010), 
        .C1(n958), .Y(n680) );
  CLKINVX1 U1087 ( .A(n1037), .Y(n1186) );
  NAND3X1 U1088 ( .A(n1193), .B(i[0]), .C(i[1]), .Y(n1037) );
  OAI222XL U1089 ( .A0(n934), .A1(n1194), .B0(n279), .B1(n1195), .C0(n287), 
        .C1(n958), .Y(n6790) );
  OAI222XL U1090 ( .A0(n935), .A1(n1194), .B0(n278), .B1(n1195), .C0(n286), 
        .C1(n958), .Y(n6780) );
  OAI222XL U1091 ( .A0(n936), .A1(n1194), .B0(n277), .B1(n1195), .C0(n285), 
        .C1(n958), .Y(n6770) );
  OAI222XL U1092 ( .A0(n937), .A1(n1194), .B0(n276), .B1(n1195), .C0(n284), 
        .C1(n958), .Y(n6760) );
  OAI222XL U1093 ( .A0(n938), .A1(n1194), .B0(n275), .B1(n1195), .C0(n283), 
        .C1(n958), .Y(n6750) );
  OAI222XL U1094 ( .A0(n939), .A1(n1194), .B0(n274), .B1(n1195), .C0(n282), 
        .C1(n957), .Y(n6740) );
  OAI222XL U1095 ( .A0(n940), .A1(n1194), .B0(n273), .B1(n1195), .C0(n281), 
        .C1(n957), .Y(n6730) );
  OAI222XL U1096 ( .A0(n944), .A1(n1194), .B0(n272), .B1(n1195), .C0(n280), 
        .C1(n957), .Y(n6720) );
  OAI222XL U1097 ( .A0(n934), .A1(n1197), .B0(n271), .B1(n1198), .C0(n279), 
        .C1(n957), .Y(n6710) );
  OAI222XL U1098 ( .A0(n935), .A1(n1197), .B0(n270), .B1(n1198), .C0(n278), 
        .C1(n957), .Y(n6700) );
  OAI222XL U1099 ( .A0(n936), .A1(n1197), .B0(n269), .B1(n1198), .C0(n277), 
        .C1(n957), .Y(n6690) );
  OAI222XL U1100 ( .A0(n937), .A1(n1197), .B0(n268), .B1(n1198), .C0(n276), 
        .C1(n957), .Y(n6680) );
  OAI222XL U1101 ( .A0(n938), .A1(n1197), .B0(n267), .B1(n1198), .C0(n275), 
        .C1(n957), .Y(n667) );
  OAI222XL U1102 ( .A0(n939), .A1(n1197), .B0(n266), .B1(n1198), .C0(n274), 
        .C1(n957), .Y(n666) );
  OAI222XL U1103 ( .A0(n940), .A1(n1197), .B0(n265), .B1(n1198), .C0(n273), 
        .C1(n957), .Y(n665) );
  OAI222XL U1104 ( .A0(n944), .A1(n1197), .B0(n264), .B1(n1198), .C0(n272), 
        .C1(n957), .Y(n664) );
  OAI222XL U1105 ( .A0(n934), .A1(n929), .B0(n263), .B1(n1200), .C0(n271), 
        .C1(n957), .Y(n663) );
  OAI222XL U1106 ( .A0(n935), .A1(n929), .B0(n262), .B1(n1200), .C0(n270), 
        .C1(n957), .Y(n662) );
  OAI222XL U1107 ( .A0(n936), .A1(n929), .B0(n261), .B1(n1200), .C0(n269), 
        .C1(n956), .Y(n661) );
  OAI222XL U1108 ( .A0(n937), .A1(n929), .B0(n260), .B1(n1200), .C0(n268), 
        .C1(n956), .Y(n660) );
  OAI222XL U1109 ( .A0(n938), .A1(n929), .B0(n259), .B1(n1200), .C0(n267), 
        .C1(n956), .Y(n659) );
  OAI222XL U1110 ( .A0(n939), .A1(n929), .B0(n258), .B1(n1200), .C0(n266), 
        .C1(n956), .Y(n658) );
  OAI222XL U1111 ( .A0(n940), .A1(n929), .B0(n257), .B1(n1200), .C0(n265), 
        .C1(n956), .Y(n657) );
  OAI222XL U1112 ( .A0(n944), .A1(n929), .B0(n256), .B1(n1200), .C0(n264), 
        .C1(n956), .Y(n656) );
  OAI222XL U1113 ( .A0(n934), .A1(n930), .B0(n255), .B1(n1202), .C0(n263), 
        .C1(n956), .Y(n655) );
  OAI222XL U1114 ( .A0(n935), .A1(n930), .B0(n254), .B1(n1202), .C0(n262), 
        .C1(n956), .Y(n654) );
  OAI222XL U1115 ( .A0(n936), .A1(n930), .B0(n253), .B1(n1202), .C0(n261), 
        .C1(n956), .Y(n653) );
  OAI222XL U1116 ( .A0(n937), .A1(n930), .B0(n252), .B1(n1202), .C0(n260), 
        .C1(n956), .Y(n652) );
  OAI222XL U1117 ( .A0(n938), .A1(n930), .B0(n251), .B1(n1202), .C0(n259), 
        .C1(n956), .Y(n651) );
  OAI222XL U1118 ( .A0(n939), .A1(n930), .B0(n250), .B1(n1202), .C0(n258), 
        .C1(n956), .Y(n650) );
  OAI222XL U1119 ( .A0(n940), .A1(n930), .B0(n249), .B1(n1202), .C0(n257), 
        .C1(n956), .Y(n649) );
  OAI222XL U1120 ( .A0(n944), .A1(n930), .B0(n248), .B1(n1202), .C0(n256), 
        .C1(n955), .Y(n648) );
  CLKINVX1 U1121 ( .A(n1038), .Y(n1196) );
  NAND3X1 U1122 ( .A(n1193), .B(n1183), .C(i[1]), .Y(n1038) );
  OAI222XL U1123 ( .A0(n934), .A1(n1203), .B0(n984), .B1(n1204), .C0(n247), 
        .C1(n955), .Y(n647) );
  OAI222XL U1124 ( .A0(n935), .A1(n1203), .B0(n985), .B1(n1204), .C0(n246), 
        .C1(n955), .Y(n646) );
  OAI222XL U1125 ( .A0(n936), .A1(n1203), .B0(n986), .B1(n1204), .C0(n245), 
        .C1(n955), .Y(n645) );
  OAI222XL U1126 ( .A0(n937), .A1(n1203), .B0(n987), .B1(n1204), .C0(n244), 
        .C1(n955), .Y(n644) );
  OAI222XL U1127 ( .A0(n938), .A1(n1203), .B0(n988), .B1(n1204), .C0(n243), 
        .C1(n955), .Y(n643) );
  OAI222XL U1128 ( .A0(n939), .A1(n1203), .B0(n989), .B1(n1204), .C0(n242), 
        .C1(n955), .Y(n642) );
  OAI222XL U1129 ( .A0(n940), .A1(n1203), .B0(n990), .B1(n1204), .C0(n241), 
        .C1(n955), .Y(n641) );
  OAI222XL U1130 ( .A0(n944), .A1(n1203), .B0(n991), .B1(n1204), .C0(n240), 
        .C1(n955), .Y(n640) );
  OAI222XL U1131 ( .A0(n934), .A1(n1206), .B0(n231), .B1(n1207), .C0(n984), 
        .C1(n955), .Y(n639) );
  OAI222XL U1132 ( .A0(n935), .A1(n1206), .B0(n230), .B1(n1207), .C0(n985), 
        .C1(n955), .Y(n638) );
  OAI222XL U1133 ( .A0(n936), .A1(n1206), .B0(n229), .B1(n1207), .C0(n986), 
        .C1(n955), .Y(n637) );
  OAI222XL U1134 ( .A0(n937), .A1(n1206), .B0(n228), .B1(n1207), .C0(n987), 
        .C1(n955), .Y(n636) );
  OAI222XL U1135 ( .A0(n938), .A1(n1206), .B0(n227), .B1(n1207), .C0(n988), 
        .C1(n954), .Y(n635) );
  OAI222XL U1136 ( .A0(n939), .A1(n1206), .B0(n226), .B1(n1207), .C0(n989), 
        .C1(n954), .Y(n634) );
  OAI222XL U1137 ( .A0(n940), .A1(n1206), .B0(n225), .B1(n1207), .C0(n990), 
        .C1(n954), .Y(n633) );
  OAI222XL U1138 ( .A0(n944), .A1(n1206), .B0(n224), .B1(n1207), .C0(n991), 
        .C1(n954), .Y(n632) );
  OAI222XL U1139 ( .A0(n934), .A1(n931), .B0(n974), .B1(n1209), .C0(n231), 
        .C1(n954), .Y(n631) );
  OAI222XL U1140 ( .A0(n935), .A1(n931), .B0(n975), .B1(n1209), .C0(n230), 
        .C1(n954), .Y(n630) );
  OAI222XL U1141 ( .A0(n936), .A1(n931), .B0(n976), .B1(n1209), .C0(n229), 
        .C1(n954), .Y(n629) );
  OAI222XL U1142 ( .A0(n937), .A1(n931), .B0(n977), .B1(n1209), .C0(n228), 
        .C1(n954), .Y(n628) );
  OAI222XL U1143 ( .A0(n938), .A1(n931), .B0(n978), .B1(n1209), .C0(n227), 
        .C1(n954), .Y(n627) );
  OAI222XL U1144 ( .A0(n939), .A1(n931), .B0(n979), .B1(n1209), .C0(n226), 
        .C1(n954), .Y(n626) );
  OAI222XL U1145 ( .A0(n940), .A1(n931), .B0(n980), .B1(n1209), .C0(n225), 
        .C1(n954), .Y(n625) );
  OAI222XL U1146 ( .A0(n944), .A1(n931), .B0(n981), .B1(n1209), .C0(n224), 
        .C1(n954), .Y(n624) );
  OAI222XL U1147 ( .A0(n934), .A1(n932), .B0(n215), .B1(n1211), .C0(n974), 
        .C1(n954), .Y(n623) );
  OAI222XL U1148 ( .A0(n935), .A1(n932), .B0(n214), .B1(n1211), .C0(n975), 
        .C1(n953), .Y(n622) );
  OAI222XL U1149 ( .A0(n936), .A1(n932), .B0(n213), .B1(n1211), .C0(n976), 
        .C1(n953), .Y(n621) );
  OAI222XL U1150 ( .A0(n937), .A1(n932), .B0(n212), .B1(n1211), .C0(n977), 
        .C1(n953), .Y(n620) );
  OAI222XL U1151 ( .A0(n938), .A1(n932), .B0(n211), .B1(n1211), .C0(n978), 
        .C1(n953), .Y(n619) );
  OAI222XL U1152 ( .A0(n939), .A1(n932), .B0(n210), .B1(n1211), .C0(n979), 
        .C1(n953), .Y(n618) );
  OAI222XL U1153 ( .A0(n940), .A1(n932), .B0(n209), .B1(n1211), .C0(n980), 
        .C1(n953), .Y(n617) );
  OAI222XL U1154 ( .A0(n944), .A1(n932), .B0(n208), .B1(n1211), .C0(n981), 
        .C1(n953), .Y(n616) );
  CLKINVX1 U1155 ( .A(n1039), .Y(n1205) );
  NAND3X1 U1156 ( .A(i[0]), .B(n1159), .C(n1193), .Y(n1039) );
  OAI222XL U1157 ( .A0(n934), .A1(n1212), .B0(n1990), .B1(n1213), .C0(n207), 
        .C1(n953), .Y(n615) );
  OAI222XL U1158 ( .A0(n935), .A1(n1212), .B0(n1980), .B1(n1213), .C0(n206), 
        .C1(n953), .Y(n614) );
  OAI222XL U1159 ( .A0(n936), .A1(n1212), .B0(n1970), .B1(n1213), .C0(n205), 
        .C1(n953), .Y(n613) );
  OAI222XL U1160 ( .A0(n937), .A1(n1212), .B0(n1960), .B1(n1213), .C0(n204), 
        .C1(n953), .Y(n612) );
  OAI222XL U1161 ( .A0(n938), .A1(n1212), .B0(n1950), .B1(n1213), .C0(n203), 
        .C1(n953), .Y(n611) );
  OAI222XL U1162 ( .A0(n939), .A1(n1212), .B0(n1940), .B1(n1213), .C0(n202), 
        .C1(n953), .Y(n610) );
  OAI222XL U1163 ( .A0(n940), .A1(n1212), .B0(n1930), .B1(n1213), .C0(n201), 
        .C1(n952), .Y(n609) );
  OAI222XL U1164 ( .A0(n944), .A1(n1212), .B0(n1920), .B1(n1213), .C0(n200), 
        .C1(n952), .Y(n608) );
  AND3X1 U1165 ( .A(n1215), .B(j[1]), .C(j[0]), .Y(n1172) );
  OAI222XL U1166 ( .A0(n934), .A1(n1216), .B0(n1910), .B1(n1217), .C0(n1990), 
        .C1(n952), .Y(n607) );
  OAI222XL U1167 ( .A0(n935), .A1(n1216), .B0(n1900), .B1(n1217), .C0(n1980), 
        .C1(n952), .Y(n606) );
  OAI222XL U1168 ( .A0(n936), .A1(n1216), .B0(n1890), .B1(n1217), .C0(n1970), 
        .C1(n952), .Y(n605) );
  OAI222XL U1169 ( .A0(n937), .A1(n1216), .B0(n1880), .B1(n1217), .C0(n1960), 
        .C1(n952), .Y(n604) );
  OAI222XL U1170 ( .A0(n938), .A1(n1216), .B0(n1870), .B1(n1217), .C0(n1950), 
        .C1(n952), .Y(n603) );
  OAI222XL U1171 ( .A0(n939), .A1(n1216), .B0(n1860), .B1(n1217), .C0(n1940), 
        .C1(n952), .Y(n602) );
  OAI222XL U1172 ( .A0(n940), .A1(n1216), .B0(n1850), .B1(n1217), .C0(n1930), 
        .C1(n952), .Y(n601) );
  OAI222XL U1173 ( .A0(n944), .A1(n1216), .B0(n1840), .B1(n1217), .C0(n1920), 
        .C1(n952), .Y(n600) );
  AND3X1 U1174 ( .A(n1215), .B(j[1]), .C(n1218), .Y(n1176) );
  OAI222XL U1175 ( .A0(n934), .A1(n933), .B0(n1830), .B1(n1220), .C0(n1910), 
        .C1(n952), .Y(n599) );
  OAI222XL U1176 ( .A0(n935), .A1(n933), .B0(n1820), .B1(n1220), .C0(n1900), 
        .C1(n952), .Y(n598) );
  OAI222XL U1177 ( .A0(n936), .A1(n933), .B0(n1810), .B1(n1220), .C0(n1890), 
        .C1(n952), .Y(n597) );
  OAI222XL U1178 ( .A0(n937), .A1(n933), .B0(n1800), .B1(n1220), .C0(n1880), 
        .C1(n970), .Y(n596) );
  OAI222XL U1179 ( .A0(n938), .A1(n933), .B0(n1790), .B1(n1220), .C0(n1870), 
        .C1(n970), .Y(n595) );
  OAI222XL U1180 ( .A0(n939), .A1(n933), .B0(n1780), .B1(n1220), .C0(n1860), 
        .C1(n793), .Y(n594) );
  OAI222XL U1181 ( .A0(n940), .A1(n933), .B0(n1770), .B1(n1220), .C0(n1850), 
        .C1(n793), .Y(n593) );
  OAI222XL U1182 ( .A0(n944), .A1(n933), .B0(n1760), .B1(n1220), .C0(n1840), 
        .C1(n793), .Y(n592) );
  OAI222XL U1183 ( .A0(n1830), .A1(n967), .B0(n934), .B1(n943), .C0(n1750), 
        .C1(n1222), .Y(n591) );
  OAI222XL U1184 ( .A0(n1820), .A1(n965), .B0(n935), .B1(n943), .C0(n1740), 
        .C1(n1222), .Y(n590) );
  OAI222XL U1185 ( .A0(n1810), .A1(n964), .B0(n936), .B1(n943), .C0(n1730), 
        .C1(n1222), .Y(n589) );
  OAI222XL U1186 ( .A0(n1800), .A1(n968), .B0(n937), .B1(n943), .C0(n1720), 
        .C1(n1222), .Y(n588) );
  OAI222XL U1187 ( .A0(n1790), .A1(n969), .B0(n938), .B1(n943), .C0(n1710), 
        .C1(n1222), .Y(n587) );
  OAI222XL U1188 ( .A0(n1780), .A1(n970), .B0(n939), .B1(n943), .C0(n1700), 
        .C1(n1222), .Y(n586) );
  OAI222XL U1189 ( .A0(n1770), .A1(n970), .B0(n940), .B1(n943), .C0(n1690), 
        .C1(n1222), .Y(n585) );
  OAI222XL U1190 ( .A0(n944), .A1(n943), .B0(n1760), .B1(n963), .C0(n1680), 
        .C1(n1222), .Y(n584) );
  CLKINVX1 U1191 ( .A(n1155), .Y(n1075) );
  CLKINVX1 U1192 ( .A(n1042), .Y(n1214) );
  NAND3X1 U1193 ( .A(n1183), .B(n1159), .C(n1193), .Y(n1042) );
  NOR2BX1 U1194 ( .AN(n1158), .B(i[2]), .Y(n1193) );
  NOR4BX1 U1195 ( .AN(n1224), .B(i[6]), .C(i[7]), .D(i[5]), .Y(n1158) );
  NOR2X1 U1196 ( .A(i[4]), .B(i[3]), .Y(n1224) );
  CLKINVX1 U1197 ( .A(i[1]), .Y(n1159) );
  NOR4BX1 U1198 ( .AN(n1225), .B(j[3]), .C(j[4]), .D(j[2]), .Y(n1215) );
  NOR3X1 U1199 ( .A(j[5]), .B(j[7]), .C(j[6]), .Y(n1225) );
  NAND3BX1 U1200 ( .AN(n1081), .B(n1153), .C(n1259), .Y(n1155) );
  CLKINVX1 U1201 ( .A(n1040), .Y(n1043) );
  NOR3X1 U1202 ( .A(n1027), .B(n1061), .C(n945), .Y(n1040) );
  CLKINVX1 U1203 ( .A(n1069), .Y(n1030) );
  AOI211X1 U1204 ( .A0(state[0]), .A1(state[1]), .B0(n1033), .C0(rst), .Y(
        n1079) );
  NOR2X1 U1205 ( .A(n1048), .B(orig_ready), .Y(n1033) );
  AND3X1 U1206 ( .A(n1259), .B(n1059), .C(n1228), .Y(n1149) );
  MXI2X1 U1207 ( .A(n1229), .B(n1230), .S0(n1058), .Y(n1228) );
  NOR4X1 U1208 ( .A(n1231), .B(row[3]), .C(row[5]), .D(row[4]), .Y(n1230) );
  NAND2X1 U1209 ( .A(n1053), .B(n1054), .Y(n1231) );
  NOR3X1 U1210 ( .A(n1232), .B(n1056), .C(n1057), .Y(n1229) );
  NAND3X1 U1211 ( .A(row[2]), .B(row[1]), .C(row[3]), .Y(n1232) );
  NAND2BX1 U1212 ( .AN(n1640), .B(n1081), .Y(n1227) );
  OAI2BB2XL U1213 ( .B0(n1248), .B1(n1233), .A0N(N2287), .A1N(n1234), .Y(n583)
         );
  OAI2BB2XL U1214 ( .B0(n1247), .B1(n1233), .A0N(N2286), .A1N(n1234), .Y(n582)
         );
  OAI2BB2XL U1215 ( .B0(n1246), .B1(n1233), .A0N(N2285), .A1N(n1234), .Y(n581)
         );
  OAI2BB2XL U1216 ( .B0(n1245), .B1(n1233), .A0N(N2284), .A1N(n1234), .Y(n580)
         );
  OAI2BB2XL U1217 ( .B0(n1244), .B1(n1233), .A0N(N2283), .A1N(n1234), .Y(n579)
         );
  OAI2BB2XL U1218 ( .B0(n1243), .B1(n1233), .A0N(N2282), .A1N(n1234), .Y(n578)
         );
  OAI2BB2XL U1219 ( .B0(n1242), .B1(n1233), .A0N(N2281), .A1N(n1234), .Y(n577)
         );
  OAI2BB2XL U1220 ( .B0(n1241), .B1(n1233), .A0N(N2280), .A1N(n1234), .Y(n576)
         );
  OAI2BB2XL U1221 ( .B0(n1240), .B1(n1233), .A0N(N2279), .A1N(n1234), .Y(n575)
         );
  OAI2BB2XL U1222 ( .B0(n1239), .B1(n1233), .A0N(N2278), .A1N(n1234), .Y(n574)
         );
  OAI2BB2XL U1223 ( .B0(n1238), .B1(n1233), .A0N(N2277), .A1N(n1234), .Y(n573)
         );
  OAI2BB2XL U1224 ( .B0(n1237), .B1(n1233), .A0N(N2276), .A1N(n1234), .Y(n572)
         );
  OAI2BB2XL U1225 ( .B0(n1236), .B1(n1233), .A0N(N2275), .A1N(n1234), .Y(n571)
         );
  OAI2BB2XL U1226 ( .B0(n1235), .B1(n1233), .A0N(N2274), .A1N(n1234), .Y(n570)
         );
  AOI21X1 U1227 ( .A0(n1069), .A1(row[7]), .B0(n1061), .Y(n1031) );
  NOR2X1 U1228 ( .A(state[0]), .B(state[1]), .Y(n1061) );
  NOR2X1 U1229 ( .A(n1065), .B(state[0]), .Y(n1069) );
endmodule

